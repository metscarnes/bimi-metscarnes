<svg xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" width="1920" zoomAndPan="magnify" viewBox="0 0 1440 809.999993" height="1080" preserveAspectRatio="xMidYMid meet" version="1.0"><defs><filter x="0%" y="0%" width="100%" height="100%" id="5d28c88027"><feColorMatrix values="0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0" color-interpolation-filters="sRGB"/></filter><filter x="0%" y="0%" width="100%" height="100%" id="c0d8f5bb04"><feColorMatrix values="0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0.2126 0.7152 0.0722 0 0" color-interpolation-filters="sRGB"/></filter><mask id="bac4022113"><g filter="url(#5d28c88027)"><g filter="url(#c0d8f5bb04)" transform="matrix(0.75, 0, 0, 0.75, 0.00000622222, 0.00002)"><image x="0" y="0" width="1920" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAB4AAAAQ4CAAAAADNuJ6fAAAAAmJLR0QA/4ePzL8AACAASURBVHic7N3XdxxHuq/piMwsb+G9B72RRFKiWqKkltTyts3pOWtuZs1fOrNmzT577XZbLU8PgAQBwgNVhfIZ5wKkSFE0MJUZmZHvc0FRbHXVJ6EyfxWREV8IAQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAIJam7AAAHIqWwhBJSuEJKoZRwhZBSCSGEUI/9Y47b1lQhgH0hgIFgiiXSuXws5sRs27HrbStr1VwnZQvbEnFRt2Nus2E5dsu1a5VU0qnUhWXJVt1OZ9bq3THRzBdKO5WUXSnXZLVUqdUaDfIYCBYCGAiKWD5tS6GEbTvxTGF4IJMvWk48FovF7EbLjclGu+3aMdsSjmhbtmy3LMtyVbxRi8dj9ZZl2ZbbshLpUjMfk7VEtlGtOKperqvd7Wp1Z2tt13Uru41YwqpVarulmu5/WyDyCGBAO9uJJ9KFgdmpgXhbtFuukHY8W8g0093KjsecuC0tt21JW7UadvJwb9GuVXZbbrVUSibE9ura2tLt5fXduquEfHzeGoCPCGBAEyvX258QdjJtx/t7evt6M+lETLhCKSWEtBzHce24kpa0LCmkUkJKoVxpKSGkUL9cuerp1/BvUrXVarvKbbuWJVy33aytLt1Z2Haa7YKsbm+urW1WXQ//VQE8BQEM+MxJJxPpTDzVNTY5lhHSSQo7nUqmk3HbEk8k597wVArxeNCq/QTwbxJYCaEe/Jm0hBSqWd0qu81mSlV3d+/PL5fK5Xq9Wt6t7TIiBvxBAAN+Sg/OzAz1Zgs98Vw2l9/7M1cJIaQlf3U9KiFVJ6/PB7GtHv+Th38um7Vqs1baLZVW1zdvXVssMxoGfEAAAz6QmWzGsuPJdP/5s8PZmBNL2E7csR/EoRJi71r09Xp8lMVSKOG2W61Wq1GrXvtmebssG6XSzs6On+UAkUMAAx6LZ4q9IzMD3SnhWvH04GBvXCkhhPzVxbeXhkG4HnfLu+UdVd1cX1tcvFferdWrTd0lAWYKwgUPGMrq6u/OZfsGhmbGuuK2EkpIy3ZsGZy0feDxiWmlVLslpFTt2t079dLGxtq9u0sbbCIGOi5A9wDAHIlcNh2LF85OjuVj8WQ2n0vYQij5cBWU3uKeZ2+NtRLCEkq0Wo16rVaen7+9UG+WtrY2GAsDHRTgOwEQSnYi2zc8O5kQDZEdGpsoxNReqkklgjf0fZ4He4Rlq7qztdFwN5cWri4slZuMhYEOCcmtAAiDZN9ILteXH57qyadjUkk7kUg6UohHm4lCSCm33Wq6ym01b/94b7O8eu/OBjuVgA4I600BCJZYPpPtOjE8lMwWcrnuVDzu/GpZc0d3FPlMPfxFNas7pfLW1au3V7bXtjVXBYRfeO8KQGBY3ccuDsXj6ZH+nkwmJYVQrmXQpfVovKuUUqqyNX9n7fpP1zdrbBcGjsKguwSggezpz6Z7T50b7pG2nUrEbceW4tn9qUJOKSGE267WquW563eW1u7dLekuCQgvM28TgC/She7jF8bysa5CsZh5eKyB0dfUgy8WSrit3c21O7d/nr+7sskTYeBQjL5ZAB7Kj5+e7MpMTI2kpZTSklJEIIDFg6fBSgq31W5Vy0s/Xb96+26JpdHAwZl+swA8IPtHuzJjF8azyVg2l3GEEDJa15JSUghXqXarWinPXb95f311ZY0nwsDBROmmAXSATGZ6jr0+XMz09fXb1mOnG0TqWlKPPehW9a27c/M3ry6scIgDcBCRumkAR2QVZmbGh/smRxKOE485D/tr6C5LL6XcVrO288Othfn5O5s0ywL2K+K3DmD/4n0jI1NTQ73FTDEvpbSEEFxB4sGT73azvr09f/Xu/aV7K2wRBvaF2wewH3Z+9Pjx6cmh3oJtW6HubNVpjx+pWNtcuDF3/ertLcbBwItxEwFeKNY7PTs9PDxayCTiMclV83RKCNVu1qr3/vHD3XvL67u66wGCjlsJ8Hy9Iz0j4yPDg8VCMWZxyTzH3sos1dpZvn1naf7W2sqm7oqAQONuAjxHov/U7PHp8aFswlJCCvngvD481V7XaKlarUZt84e569durNV01wQEF7cS4Fmy48enxsYGevPplGPLSHTZOLq9Ph1uq1mrlL795t723CJrsoCn434CPI1d6B6YOT4+MtSXSUgpRETaXHXAozbYbntl4dbV23ML6xWdBQFBxf0E+K34+PHZmenRvpzj2HLvWEFDj1fwlHJdt7Jw9fq1G7fWW7qLAQKHmwrwBHtoZPrU1HBfVzblsOrqCB5sEK7s3P3HtXtLiys0jAZ+hZsL8CvZ/vGzMzMTQ7n43sgXh6WEEEpIqZS7c3v+zrXv5lZZkgU8hvsL8Ei8f/rczMxQby4Vty3dxRhDCbfVqK/81w93526v6C4GCA4CGHioZ2zixPT4UH826UiujM5Sql3d+OmfP/ywtVXSXQsQENxmACGEELHi8PljJ6bH8gmGvl5R6//xn/W1W7c36rorAYKAAAaEkIPHpk5ODvUVMinH4qLwjFsvN+/98MONufkN3aUA+nGvAXL9QxdmJ0cHcynC12tKtKqrP/7r5o27KwyDEXXcbxBxVnby2MkzxyYf9dvgovCYaldu/vuna1cXOK8B0ca9BpHWPTVxbHJkqDufs21J+PpEufXdlX9+Oz8/t6p01wLow/0G0eUMDJ2fnZoYKWYedrvigvCNqi1999MPP9/acnVXAujC/QZRlZw4d/r41Gg2GbMsJSQXg8+U29z5+99u3bl5v6m7FEAP7jmIpv7pkycnx/q68g8abnAl+E+1GxuLP/5w/Q5rohFN3HYQQXbv+MWTx6f68pYl1d68M1eC/5SQ7WZ96+o3334/x5mFiCBuO4ic2PjLJ47NDnSnHMui45VeSrmtRuXv/3H3zo37PAxG1HD7QbTYgyMDl6ZHh/rTcakU+RsE7Xrp1n9/f/PWQkN3JYCvuP8gSqyeM2dOn5gYSDgWK54DQynZqt759se//7xEBCNKuAchOhITp04fnxjOZ1NMPQeKkm67Ud785u+3b81v6S4G8A23IURFcmTm1dnp0e6spOFk8CjhNivrP/7rx++XWY+FqOBOhGiIjZ9/9fTxvrxN+gaTUkq1m5Xv/p+FO9dYj4Vo4GaEKMjNnD91bGygKxkTfOgDSgmhlNus/PzND9duLLV0lwN4j3sRzJceOPH2ianRXEIqIfjQB5kSolX54V83v7+6wnosGI97EUznHD/90sXp7kzcshSf+GBTQgi33aps/eNfP/y8SATDcLbuAgBPpSbPvf/JpenBbNym4VUoSMtJpIcnkvm80yCCYTTuRzBZbODcxYvHhzKO5LiFcGmVfvxp7rvvl6q6CwG8wx0J5kpPz5x8+WRfbm/bL5/18FBCufVq6e//uH7jLhuDYSxuSjBVcmLmyrHp/kLStpTgox4qSgghhFtZ/Pbbqzdv7WiuBvAIdyWYyRp8+c1zx/rzllDs/A0t1br7zX9/+9/LPAuGkViEBSMNvvbFhxdmezOOlHSdDCslhEiNHO9LF1SJ1hwwEAEMA+VPvP7p5fNjvUnyN+ycZG70WDEj6ru6KwE6jgCGcWLjb//h0wuzXQnmnsNNSimFtJM9k5PZvCo3ddcDdBgBDMM4Mxffv3JxtjftEL8GkFJK28lPddvFdJs9STAL9ygYRfYfe+ns6cnetO5C0FGqtvDtTzd/ml/jWTAMQgDDJIMnT585NdaXiFl8tk2ilNuulu79/ftrP3NSEszBFDTM0Xvxtd+9en66N+PQd8M00omlu2eHszmnwXIsmIIAhimSU6/+7sqbp8eyjhKS/DWKFFJYdjw7eqonnm2X2rrrATqCAIYZ7Nk3f//7V0/0px0p2XtkHPlAYni0mukuV3TXA3QCAQwj9J1/43eXzo/3JG3i12DSindN9HfH1C57kmAAAhgGSBx78713Xz/el7AIX7MpIXOjJ3LpQnOXeWiEHncrhF5q9uTZ05Mj+YTN59l8SqlWaePW37/77hYdohFyjIARcsnRS++8efncWHfcEnyjNJ8UlpMujp3IOe0t5qERbo7uAoCjsKZOnT97qr8Qt11WPkeDFEJYyYEPsq5cYFMwQo0RMMKs5/U3r1w8OZpP2JL8jRQrPthfSMTrdKdEiBHACK/Y1FtX3nhtZiBtCzpvRIkSQojY8Ewm092sMQ+N0OKmhdAae+nc+eODhZjD4DeClBJubf2b///mwo1t3bUAh8MIGCHVdeq9K5dOjxYTNvkbRVJYVjw3OV7Ippolpbsa4DAIYISSNfmHj9994/jAXuMN3dVAAymEsGL9U73JbLvCjiSEEQGMMBp5/ct3X54qxsneSFNCiFj/RK+TETush0b4sA0J4ZM79vprx6YKSYuZR1jxgUJuoD9/Y0t3JcBBMQJG2Mjpj7768KWpYozGG1G3d0CDFRuZTKaSNKdE6BDACJmhV9797NxEMWFLIZiBhhBSWqmxnJuMcVIwQoYARqjEjr/7l3fPjORjllAMf/GAnRgbKiYz7TKDYIQJAYwwGb384duXx7KOFILFz3iMKh6fLSinxiAYIUIAIzwyJ1/5y7vnupK2xcNfPMGy08P9yaRdq+uuBNgvAhihMfDax5+8MZZ1JFt/8QS59yR4NNZll6ssjkdIEMAIieTLn3/+1plc3CJ98VtSSmnZuWNdIp3ihAaEBAGMcOi//Ne3zo7kHfIXzyCldJKjQwkr7tKbEqFAACMM7DN/+Oubp7uThC+eRwm7d7LZHGyWWrpLAV6MAEYIDP/u91+d7U1ZxC+eS0ol4jMnhmOyWtFdC/BCBDACzz7+ztfvn+gjf7EvTn4kayWadIdG4BHACLripbc+fWsoy0cV+7DXm3Jo1HbcMkckIeC4qyHY5LFLV/54qjtusfMX+yOlZed7m1asxjQ0go0ARqDFT3/w2YdTXY6k9Qb2T9rdA8lYolliGhpBRgAjyHovvPvphcGExbkLOAglRHZiMpdVuzXdpQDPRgAjuJyplz/+/FhXks6TOBgphHS6RgvJeJUtwQguAhiBlX7lrbc+m846kuEvDkhKIWVmfNxxWluckISgIoARUHL6jU8+fa0nbpG+OAQphbQy2d2W4ngGBBUBjGBKnfjdV29OdSfIXxySlDLWPeTEHZpyIKAIYATS4KUrn747kLHp/IzDU8IqTPa0rWaZ1dAIIgIYAZQ69dZnn53IxSzdhSDUpBTS6RvLxUWV1dAIIAIYwVN85ZPP3hrKMfuMo5JC2N1D6bjc3WU1NAKHAEbgTLzxxefHu2LkL45OWpaVHut3ks0dVkMjaAhgBEzy9Ht/vjycc0hfdISUVqyrxxKNbRIYAePoLgD4lfxL7/1hqp/4RedIO3OqYNvqJg+CESyMgBEok29++slMIU7+opOUzPQ7datW1V0I8DgCGAHiTF3+y+9H8jHyFx0lhZXpy2fTdU5nQJAQwAiO7NlTX33RkxK0fkaHSaHS01M5p7nT1F0K8AsCGIExdemj/+ti2hY030DHSWnZyeFkMtPgdAYEBgGMgEie/uDL30/mbcnwFx6Q0oqnxwqO1Sq3dNcC7CGAEQz5y3/56NxYkt6T8I4VHxqsJzIl1mIhGAhgBEL/Sx+/O9mVIHzhJSkL410Zp7qjuxBACAIYwTB68bPPZgtx3WXAcEpY+dGCcBoVpqERAAQw9JMzZz//U1/SYvUzvCWllFZPfzquyjTlgH4EMLRLnn7rT+/3Jchf+MGyc72usttlVkNDNwIYuhVe/fijN/oci+VX8IV08mOWSrVL9IaGZgQw9JIzVz7+8EzW5uhf+EYmJ0ZaCavU0F0IIo4AhlaJ02//6fXRos3oFz6SsZ6uWMKtsB8JWhHA0Cnz8pdfXhjMSB7/wk9KyO4xyxHbu7orQaQRwNBo5LXPPpooxIRgAAw/SSlkoi9pyQZLsaARAQxtkqff/uPbU4UY41/4TgorM5BSbr3M+UjQxtFdACIrf/mDK2O9cQa/0EEKkb2Ua4rkHNPQ0IURMDQZuPzVG9PFpEX+QhPp9BYcW1XqugtBVBHA0GPk9a/en+yKEb/QRglroF/F5C5jYOhBAEOLiYuffdqb4ukvNJJSiOxUd1rtcjgDtCCAocPU5T++35ewyV/oJa1EV7wp6iUWQ0MDAhj+k8cu/+WDbsdi9xH0klJaqeFMM93YoS8l/EcAw3ex0+/936/kHHo/IxCsvoGYUPSlhP8IYPgt9fIHf53qiVnkLwJBOsVeK96sshQLfiOA4bOu17/89EQhxvgXAaGEzI731K1GSXcliBoCGP6auPzx2+M5m/RFUEgpZLyQkTG129RdC6KFAIaf7GNXPn9/tOiw/BkBIqWVGkxYSVWiJwf8RADDR8659z+9PBRn+TMCJzbQJ2y7xAGF8BEBDP/Ez77z5dmeJPmLAHK6uhzpViq660CEEMDwTeLsHz67UExI1l8heJSQhaJrq03GwPANAQy/pF567+uTOccifxFAUgqZHkjGVIXF0PALAQyfZF/95KvZfIzTjxBQUshkj+OoCp2h4RMCGP7IvPrnj2YyDqNfBJaUMtmXV62dsu5KEBEEMHyRfuXdj0ayNvmLIJPCKcZst77D2QzwAwEMP2TPvff5iVyM/EXAWfHeRFvWt0lg+IAAhg/yL1354nTKpvsGAk5KGesrtuUuCQwfEMDwXv53n38+xfNfhIK0u2LCrW2RwPAcAQzPpV768qPptMP6Z4SCdHrSSpW3dNcB8xHA8Frm/LvkL0JE2T0D1m5lW3cdMB4BDI9lXv7w65Np1j8jPKTMW5a7u6m7DpiOAIa3si+/95czSYv1VwgNKaTV3dVolOmJBW8RwPBU7tWv/+dIUpK/CBEphZ0XymqwEgueIoDhpdyrn342lLZ0lwEcjJROtxNr8RwYniKA4aHUxQ//PMb4F2EUH+jdqjXLru46YDACGN5Jnv/9n4dTFuuvEEZWoVgU9U0SGJ4hgOGZ9Cvv/vlMkvXPCCUlrb6uZrPMc2B4hgCGV7KXPvw/j8V5/otwklLKTLpeq5cYA8MjBDA80n3p878Mp8hfhJe0Cpm8qm2RwPAGAQxvjL356dejCaafEWJK2H19rUZ5hwSGJwhgeME5894fP+iJk78IMymllYm3mw0SGJ4ggOGB2PlPv7jUxfgXYSel1RWLtWvbJDA8QADDA+c+++x8D8cPwgDS6RvcbVU4HxgeIIDReWOvf/5ShtOPYAYrG7cqtR0SGB1HAKPjht//8vUi239hCGkX4sKqsh8YHUcAo9N63v+fr/VYkgCGIZTTNyIaW/SFRqcRwOiwzKWvrhTj5C+MIYWVrNXr5bLuQmAaAhidlbr08RfD5C9MImUsUW81tqu6C4FhCGB0VOL8e/9jJMb5RzBMKt2y3Y267jJgFgIYnZQ48/4fZxMW+QvDWOmCELsbTd11wCgEMDooff7NP11g/hkGsosp0SyvshQaHUQAo3MyFz79P44nOP8XRsoXKvWtLd1VwCQEMDomc+HTLyfTFh04YCQr4dZrOyyFRucQwOiUzMUvvppO2uQvDOV0O7uNnV3dZcAcBDA6JPnyB5+Mp2iABXPFsrFqfaOhuwwYgwBGZ8TPfvDh+TT5C5MlC416ebOtuwyYggBGRzgn3/7qQpL9vzCaTGZb21XOJkSHEMDoBOvsh5+8kmL/L0yXiceaO5u6q4AhCGB0gHXqDx9fzrD/CMaz8+lmZYOFWOgIAhhHJ89//P6lHPkL40lhFWVre5OelOgEAhhHd/Ljj1/Js/4KESClk25vV7ZauguBCQhgHNn455++mnPIX0SBlKmu7Vpli4VYODoCGEfV/9an54vkL6JCJrsb9d1tukLjyAhgHFHy8mfv9CTIX0SGVczIWpmu0DgyR3cBCDn77LtX+uPsP0KEyBOF3d3dFd1lIPQYAeNoTnz80XSKBhyIllQ6VStxLgOOiADGkYy88eXpLksQwIgQJWXR3t3drOkuBCFHAOMoim9+9VYhRv4iUqSUsUSrVN1kMxKOhADGEWRe/fTKYIwJaESNlKncdr22yWYkHAUBjMOT5754byxNByxEkMyLuqrQFRpHwSpoHN7oq7/rT+kuAtBCnXaS1Z37ustAmDECxqH1vPnF6S52ACOi7LSs0RUaR0EA47Byl/708lhCEsCIqHh3o1LaaeouA+FFAOOQMq9+9sZQyrLIX0SSFDIhm+36Rlt3JQgtAhiHk7zw0QcTOYf8RVRJKTOJZqO0RVdoHBIBjEOJvfTxlzMZxyZ/EWFOIVWqlkq6y0BYEcA4DPnKJ1+P5DgCGBFn51q1VqmiuwyEFAGMwzjx+afHOQIYkSfjedWsrrEQC4dCAOMQZv704Wye/AVUsk/V1zd4DIzDIIBxcH1vf3KiN876K0DIZLKxVtnWXQZCiQDGgTlXPr3Sl2L8CwghZDGx3KyxEAuHQADjwM588NFonPwFhJBSynij2irv6q4EIUQA46DG3/9qNkv+Ag8kinVV26EnJQ6MAMYB9b/59eU8BxACD8lcwd4t0xELB0YA42By7//l7axD/gKPZFK7u9tbuqtA6BDAOJDYpa/eGSJ/gcdZWWttc72huwyEjaW7AITLqU/f6mf/EfBrzujAQB93UxwQI2AcxODHX0yn+dAAv6bidrqyxV4kHIyjuwCESebyH6azjmIEDPyafSpzf2WdldA4EAYz2L/YxS/eHKQDJfAb0kqVyiusw8KBEMDYvzOffDySIX6BJ0lh2WqrXCrrLgShQgBj36b+8PGFNPkL/JaUdq5VrpWqugtBmBDA2K+Bj756KStpwQE8lZNrb5R3WrrLQIgQwNin5OWvL/Q5BDDwdDLdtVGtbru660B4EMDYpzOffdifkqzAAp5BZq1ajb1I2D+2IWF/hq5c7kuSvsBzHK80trYruqtAaDACxr5kXv3j6QGbAAaeSSkn197Z2GISGvtEAGNfXvrT7wYT5C/wbFIoJ7dbWmMvEvaJAMZ+DL370WSODwvwXNJKlUrbG03ddSAkuKdiH1K/++RyMaa7CiDYpLScZHm7tKl0V4JwIIDxYvb5z98Zjkl6QAMvko6t7ZZYCY19IYDxYjMf/nEkK9kCDLyQlRW7lU1OZcB+EMB4of63/no2JwX5C7yQsvsbO1vbbd11IAwIYLxI8eP/cb7g0IID2Bc7myhvbuquAmFAAONFLvzlwnCc9AX2QwqRSq1trDV0F4IQIIDxAuN/+HiUMwiBfZKW7Wxs72zSjgMvRADj+dK//+pcho6lwL7JRHprtcxKaLwQAYznO/fl60MOO5CA/ZMFtVIu1XSXgcAjgPFcg+99OcoZSMDB5KzyzgaT0HgBAhjPk3rjTye7HOIXOBArV9ld29FdBYKOAMZzWOf/+G5vkvEvcEAZt7myzSQ0no8AxnMc++M7kwmLAAYORsp0c6u6zakMeC4CGM/W/d4XMz02LSiBg5FCJrONWoW9SHguAhjPduHr1/rjrMACDkpKmRmo7myyFwnPQwDjmUbf+WgkZemuAginzPZGbaequwoEGQGMZ8le+ehilhXQwKFIGW/WSmtMQuPZCGA8gzz32ZuDMR4AA4ejUl2NynJZdxkIMAIYzzDy7mfDWVZAA4eWcOtb20xC45kIYDxd7PU/nS3ELfIXOCRp5Rvl0kZLdx0ILAIYTzfx1eXhpE3+AockpYxlGrulDaW7EgQVAYynyr39yUzBZgIaODxpJbvWyqtMQuMZCGA81dk/nR+OswILOBI7X1vf2mjrLgMBRQDjaYY+eX8kZ5O/wBGpra2dbd1FIKAIYDxF4rXPzxcT5C9wVPF2s7LFJDSeytFdAILoxNun+2nBARxd8rTc3SzXdZeBQGIEjN8auvLFRJ4FWMDRyVi+XFpjEhpPQwDjNxKvfvFyb5z8BY5MCjtpba9tcTQwnoIAxm+89Od3+5KsgAY6QEqZL69tb9ATGr9FAONJg1c+mE07zEADnWHJ5d3Sju4qEEAEMJ6QufjZhQFacACdIhP1nepaQ3cZCB4CGE84/v4ng0nyF+gYp7te3qAjJX6DAMavZd/4+kSOHtBAxyiRtJtbmxxMiCexDxi/dvzy6RyfCqCDpJpt37u/xrFIeIKluwAES+/FV4tMiwAdJIVl943NjuuuA4HDvRaPs859cr6fCWigk6S0nHqptE4/LPwaAYzHjbz10Via/AU6zMnvbq+v664CAcMUNB5jHXt1IqlYrQl0WtfM6FSP7iIQMAQwHtN76lwxrrsIwESjp2bGdNeAgGEKGo+krvz1ZNFiDzDQcSqZL2+v7OouA4FCAOOR419eHI1b5C/QcVIkauWtVbYi4TEEMH5RfOOrmQLxC3hBOpn65uqW7jIQJDwDxi/OvjOVIX8Bj3TPjI2wxAKPIYDxUNfFU/0J3UUAxrLGZke6dReBICGA8dDE5YmUzRYkwCvZY2ND3HLxCJ8GPDD4zmSXZAU04Bk5MjuR1V0EAoQAxh777NnhjO4iAIMpmRuf7dNdBQKEVdDYM/bRFZpQAp6yndq9NTpC4yFGwBBCCBF75dxoUncRgMmktIdnZ0e56eIhPgsQQggxemW2LyZYggV4R1qp0yemC7rLQGAwBQ0hhEi88+E0TSgBj0k7tr5z39VdBgKCETCEEGLmlYkC+Qt4zZk5NtuvuwgEBQEMIUTilVNDGUH+Ah6ThZnZ0ZTuKhAQju4CEARTr0wmOIQB8MHp+urmdd1FIBgYAUOI5KXZwRgT0ID3ZPHsiSk6QkMIQQBDCCHGLo7nLcUSaMBr0nL6TvEUGHsIYIjcpZf74nShBPwg7ZmJWRpSQggCGEKI029MFx3iF/CFHJ4+xhAYQhDAECLz2rGepMUaLMAXMj41O07fdQgacUCIPG1BzQAAIABJREFUc5+dHbSJX8AfSiTkxvqa7jIQAIyAI69weXaA4S/gn8JL56bZCwwCGOLEy4MpwRJowCdS2t39I926y0AAEMBRlzp+vCsu6IIF+EVa9uzwaEJ3GdCPAI66qYszeZstSICfxsfHWAgNAjjqkmfPFh3mnwE/qfTZk+MMgUEAR9zka6MZlsID/rImzk536S4C2nHvjbbM+1+PZ1gDDfhL2emNZc4FjjxGwNE29kof2yEAn0krNjQz26u7DOhGAEeaM/1KMcYeJMBn0klNzw5zGmzUEcCRNnFhPG0p9iABPpPO0OAYQ+Co4xlwlMXf//x4kj1IgP9krL21cU93FdCLAI6y2T+fG7E5hxDwn7Jy1c2Fqu4yoBUBHGG5Kx9O5C3yF/CfFHZ86z4LoaONZ8ARdvy1yQL5C2ghnZGxSfYCRxsBHF3xV04NsAcJ0EPameFhlmFFG1PQ0TX7+csDDuNfQA8lU7WV9V3dZUAjRsCRlb50bJD8BbRRufOnJrgEo4wAjqzxS8NZenAAukgZGzs1m9NdBjQigKMqduJ4tyPpwQHoIq300MSE7iqgEQEcVSOvTucs8hfQx3KOTdEROsoI4IiyL0z3JchfQCc5dGJ0iKswulgFHVGDX16YcDiHENDKSpbXVmiHFVmMgCPq5NmxBGugAa2UKr52ZkR3FdCGAI6mngujed01AFEnpTN8bDqruwzoQgBH0/jL/TTBAnSTdnZghGVYkUUAR1Li+Jm8xRZgQDcrlukaTuiuApqwCCuSjv3ltVyMNdCAfunK9uq27iKgByPgKLLOznTHiV8gAPpeOjmmuwZoQgBHUfe54RhNsIAAkGJ4Zox+lBFFAEfR7PkejgEGgiE5OjyguwboQQBHUO/5YwVOYQCCwR4fGmMZVjQRwBE0/WYxwQAYCAaZHxoq6C4CWhDA0RM/NpVl9TsQFPbkMeago4kAjp7Ji2NJzkECgkEJOXVmjCFwJBHAkZN65WyXwxosIChkcmqGIXAkEcCR03dxOMOPHQgIKa3kyOigo7sOaMCdOHJ6j/fYjH+BoJBWoljszuguAxoQwFGTP3M6S/4CwSGt2KnJUd1VQAMCOGrGL/clddcA4HH2iWPTLMOKIAI4Yuyxk0l+6ECgyO7jk326i4D/uBdHTM/JUYcfOhAoyh4Z74/prgK+414cMTMvDdKEAwiantGBvO4a4DsCOFoypy+mdNcA4Em5YzNDumuA7wjgaOk/081EFxA4zuD4CCcyRA4BHCly/EyOJlhAwEhp5QZGmIOOHAI4UnrPneNbNhA8Mjk5McjtOGr4iUfK2NleZqCBwFHCGhsfL+ouAz4jgKMkNniMJdBA8EhpFUenenWXAZ8RwFEy+NIJHgADASRlfHJyOK67DPiLAI6Q2Mm3u4RQussA8BvSHpoa6dZdBfxFAEfI0Mun4kowBgaCyBntYRlWxPDzjpC+2ZzNJiQgmKyx8RHa5EQLARwdsjieJH+BYFKiMDuQ1l0FfMWi2OgYePXLbn7eQFBZRbu0vqu7CviIEXB0TJwbslmBBQSU5Qy9/PKU7irgJwI4MpJjZ+KSNdBAMEkpZd/MeFJ3HfARARwZxdlRS7AGGgiu7PAIZyJFCQEcGQMni6QvEGSxqZEpmsVGCAEcFfHJYxyEBASaNTA+26O7CPiHAI6KgQtTCckMNBBkiRkaQkcJARwV4y9nHUbAQJCp9vBYj6O7CviGAI4Iu2+M6xoINCVEZmo0p7sM+IYAjojCRD+LO4CAs+J94wO6i4BvCOCImD7XbbMJGAg0KZ38+KjuKuAbAjgixs7GeAAMBJoUll3oHcjorgN+IYCjITvUxUFIQMBJaTnjQ126y4BfCOBo6J/OS9pgAUGnxMjgJMs1ooIAjgR76iznnAHBp0T37Gy37irgEwI4EnqPnaLHOxB4Sgjn2Gy/7jLgEwI4EnqneizWQANBJ6Vl5U+OxXXXAX8QwJHQdyrGTxoIPimtVP9AUXcZ8Ae35ShIjpywpWIJFhB4UqYG+jmTMCII4CgYOjlI+gLhEOubGGPJRjQQwBGQmDqTIoCBcLCzU6MJ3UXAFwRwBBTGJzmIAQiN4eGU7hLgCwI4AnK9vVLSBwsIAyVkf3+f7irgCwI4AnL9HHAGhIUS6Z6BrO4q4AcC2HxOcYwnSkBYSBkbGKMZViQQwObrHj3BI2AgJKSUTv9or+4y4AcC2HzDM5MWXbCAkJCW3TPcy0akKCCAjeeMnsxJ+lACoSGTfUUeAkcBAWy89PAJixXQQIg4Y33MQUcBAWy8wuCwxSYkIDSUsAYGBzmQIQIIYOONn8zoLgHA/kkluk6Od+kuA94jgE2XG+UoYCBUpOWMj/XorgLeI4BNVxge5IcMhIm0YoPjw2ndZcBz3JtN1zvOsyQgXCw71zU+oLsKeI4ANt3gbIw9SEC4WKmx6VHdRcBzBLDhkrMnHZZAAyFjjUwMx3QXAa8RwIbr6SvYumsAcDBK5IZ6eHhkPALYcKM9aQIYCBflKqtY5BAz4xHAZnMGh2LMQAMhIy1n9PiI7irgNQLYbOnhUzb5C4SLlJaT7JmkhY7pCGCzZae7BYuggZCRtpOMjxZ0lwGPEcBm6zud0l0CgIOTTn9/UXcR8BgBbDR7eDTBDDQQOkpYA31dXLyGI4CNVugvOFzDQPgole3qZR204Qhgo3UNd0khiGAgbKSI9/RyIIPhCGCj9c7Ygl1IQOhIKVRPf7/uMuAtAthoqW7FEmggnPrHe2mGZTYC2GRO7xRtsIBQkjLe1UU7aLMRwCZLzUw4kiEwEEaW05NnBGw2AthkI0MZfsBAOFnx7jQ7gc3G/dlg8clZjiIEQko6vd1DDIGNRgAbLDM2IyWbkIBwksWRCTYiGY0ANliykFLkLxBKUsrU5OyA7jLgJQLYYOn+pCJ/gXCS0hqZ6OUWbTJ+ugbrP53mJCQgrKTMdGUd3VXAQwSwueJDE6zgAEJLifxQL2cCm4wANlfPyFCMGWggtGR8eLBbdxHwEAFsrqHJomQXEhBWUtqJ4ojuKuAhAthcfWM2+QuEWbZnMKW7BniHADZWrGuQFVhAqKUGh9K6a4B3CGBjWbFejkICwky5A32MgA1GABsrkS+Qv0C49XcTwAYjgI3VNVMQDIGB8HKVzI12cZM2Fz9bY42dYBcwEGZSWrHscFZ3GfAMAWyqzOS0TSNoIMSkJWPdY5zHYC4C2FTdJ5LSYhsSEGZSFif6dBcBzxDApipOJRgAA2GXHenXXQI8QwCbKjsQc3XXAOBoVGyAA5HMxY/WVH3DDmuggXBTwu7P27qrgFcIYEPFuvKcYwaEnbRzqZjuIuAVAthQ6WKa781AyEnLtuO04jAWAWyoocmEzRosIOxsJz2kuwZ4hQA21MiIYxHAQMhJmS5OJXVXAY8QwGay+rssiwQGQi8xOkovLFMRwGaKdedZAg2En9vu7c/oLgIeIYDN5HTlCGAg9JRqdfcQwKYigM0Uz6YV24CB0FMq3d/NfdpQ/GDNlEyleQAMhJ4SMt7dn9ddBrxBAJup0JtkCRYQfspODo5wHoOhCGAj2YPdMZujkICwk3Ysnpsc1V0GvEG7QiMVJ6cc8hcIPWlZIj866rR0FwIvMAI2UveJLilZhAWEnpTCHumjr6yZCGAjZQdiQnEcMBB+SllD3QSwmQhgI+UHbaHIXyD0lBJWOkMAm4kANtLYhM34FzCAFNK2nbjuMuAJAthEVk+CTUiAEaRlW1aX7irgCQLYRDIZt1gEDXTCw5ZyuhY1Sttx5BBz0EYigE3kbCf4wQIdIR98l5VSCaG0dHhNZkeL/r8rvMd92kSpqsv4FzCF7BpiDtpIBLCJ8rIpBLuAgY6SQs/SRuUW+gs63hheI4BNNPh2LyNgwAN7F5av89BKiaG+PE0LTUQAGyjed9whgIFOU2ovgf2eXZKpbJJVWCYigA2U7O+xJaugAS/4PgaWlpNSTsy394N/CGADpYpF4hfouMcvKx+vMGkl8tm0f+8H3xDABsqNpchfwBtKiF9HsfdkrC+f9/MN4RMC2EDDF5MsgQa8sXfMmM9XWDLLMmgTEcDmiXeNsGAD8JD0dz+SEoXhHh4CG4gANk8qnbK09c0DDKf8X+DoupkxAthEBLB5MoM53SUAxnqYvn5+xbUsm3UdJiKAzdM1FBOaWvYA6DxpJVIJrmgD0V7FPMMjllB8swK8o3x9CmxJmU9ySRuIADZPs8XwF/CUz1eYcotJ7tUG4luVeWouE9CA53xc6KjcbDru27vBNwSweRI9Ws4sBaLFv8XQrtvODrO00kAEsHGs0RHGv4BJlIoV+pmDNg8BbJzE2AABDBhESssuDmd1l4GOI4CNE7djBDBgEjvuJEZoRmkeZjWMk8ulOAsJMIiUQhX6eAhsHgLYON1DCYsABoxiZbo4D8k8TEEbJ8UeJMAXPu5DEvlepqDNQwCbxsrQNBYwi1LCyaV0V4GOYwraNKmeYd0lANHg21ddKYQd45BR8zACNo2T4tgywDBSOnGbqS3jEMDGkQ7XKeAT35rO2ZzGYCB+pqZplfw/LxyIKt8uNovNDQYigE2THynQCRowjBK+HoAIfxDAphl+u0D+AqZRTGwZiAA2TXaERViAWZRSsq+bK9s4BLBp4ikeFQGGUUIm8pzGYBwC2Dh1H7cnAnjAyyc/UkpLZno9fAdoQQCbptViBAz4z9PLTkohnX4v3wE6EMCmcZLs1weMI2OZnrjuItBhBLBhEiMjtBcFTKNUvL8nqbsKdBgBbJh0lv36gHmUyOUTuotAhxHAhknE2QUMmEepTI7JLdMQwKbZXHV1lwBEjedfe5UQvWwENg4BbJhEPq27BCByPH/sI4WIMQA2DgFsmO7povffxgE8hbdbgVuNtoevDx0IYMOMHEuyBgvQwtNLT+VsL18eOhDAhukasGiEBRhHKR+eNMNnBLBhLE4DBkzkttsEsGkIYMPYbEMCzKNc1x5M6a4CHUYAm0U6NgEMmMjJscPBNASwWWTaFooIBgwjLTtWyuuuAh1GAJtF1ao8AgbMI23H6snorgKdRQCbRW1VdZcAoPOkHc/2FXRXgc4igA1TqbIMGtDFs8c/UgoRy+a8ennoQQAbJlEgfwFdPLz4lCp28RDYMASwWezuXtZgAeZRbTXAM2DTEMBmiQ1YLgEMmEdKZXEcg2EIYLPYKaloWAcYR1qWY3G/Ngw/UMM0SF/ARFLGbRZ4GIYANkvzbs3iIgUMpFjeYRwC2CxqpWWRv4AGSglPDyxymy1OOjMMD/XNkjrXo7sEIJq8DUel2i0mt0zDCNgs8b44q6ABAyklHe7XhmEEbJZ43G0LJqEBLZSHw2AlrBT3a8PwjcosmbTLCBjQRErvelHaTqzJtW0YAtgsKUvxnAgwkLQcNgKbhikNs1jbIk4AA/5TUggvV2IpYSVsz14dWvCFyih2cSRB/gIaeH7htRu1NnPQZiGAjZIs9iV01wCg85RqNRpt3VWgswhgo8RzfTbfkQEDuc1akqvbMASwUZw4W5AAI0kp6m0ub7OwCMsoUtpcoYCBpGU7u03dVaCzGAEbRcmY7hIAeELaKYfv12YhgI1iWS1Xdw0AvMFxSKYhgI1iO80W1yigjXdnBkq3Xa5ydZuFADaK23ZYhQXo49nlp9xmPc4UtGEIYKMoEeMnCmjkWUS6bivOEg/DcLs2ipWgEzSglYdXIAFsGgLYKJYjWacBaOTZ9Wc5iVqT79dmIYCNYjuslAT0UEoIobxKYCmduOtywzYLjTiMolqK71SAFp6PTu3+LCNgs3C3NkqbTUiAXt6tgxb9RQLYLASwUVzacABaeReRrirkuWGbhZ+nUTx7AAVgH7y7/pTbbjddRsBmIYCNkshZrMECNPLs+lPSiSXjXr06tGARllGKQ7ZS3i8GAfBUUgnl0fUnE0p05ze8eXHoQQAbxW1KSSsOQBclPWsFbcVt18579OrQgyloo7hKkL+AFsrbJRjSScQTedvDd4DvCGCjxJLEL6CBEkJKJaWn34CtdIpmlEYhgI3i1lmCBWjgxzdf1WjZ3LGNwjNgo7RrLgkMaCL3RsKevX6j5dlLQwsC2CiWLZRXizABvJCHV59SqZx3rw4dmNAwimWzBgswlmSGyyyMgI2iLHYhARp5OAUtRatBAJuFADYL88+A556bsl5OQjcJYLMwBW0UpqABnTzOx1ab41aMQgAbxXbIX3RW5IdcT+mu/qwHPUp5ex6K3Wy1vXt1+I8paLNIWkGjsyL/cTrYfwAv/3OpVq3CCNgojIDNYnMYEuAF9Yzf/4qnayCVqjdK3r08NCCAjeIkPesFj4jiA7VH/vb3j/2nUQ//3MsDgVtWrOzZy0MHAtgozSozhoBP5FN/65322lbVj/eBbwhgo1RLnIYEaPHLINgjUqrV5bpnLw8dCGCjtF1GwOgsPlD79GD+2btvwNLuSXn12tCDADZKu84iLMBQ0hYsgjYLAWwUxWlIgB+e+k3X00VYQrm1Npe3WQhgoyTyigQGOu43V9WzWnF4NgGtXCUKBa5usxDARomnhWISGvCFz1eaEvE4F7dZCGCjWEqyDBrosAeHbD9Mv4d/fcqV5t0ktJSWKLMLyTC0ojRKo6zIX6DD9q6pX6aXn3mJKS8fAkshXTpBG4YRsFFqJX6iQAc9eqKzv8e7Xs4RE8DGYQRsFGVZDICBjnksT597ZSkhhBRSCS97wbpbdKI0DAFsFMsmfwFtPD0LSal00sPXhwYEsFGsmJcbIYCo2e/FJJ/yu85SypW9bEMyDE8MjWIL+fQOAQCO5rnXldrXP3UUUgpV5xmwYQhgoyi3wTYkwEhSuHy7NgwBbJTWbo38Rcdx3xcvmFt+sP9IefoASLLEwzQ8AzZKo843KnQe9/19kkJ59h9LSrnb8Oi1oQn3a6Mot6W7BCDaPOzEUSWADUMAGyWey3m5DxHAs8jHfvWGarEIyzAEsFEUx5UBplKNpu4S0FkEsFEalSbbgAETKekSwKYhgI3SKK3rLgEIvwNNJKnHNwF7NwWllKrxDNgwBLBRGtUac9CAr3za+SdFe7fuyzvBN2xDMkqj1lSKXSPA0TzjCnrRHiP57P/r0UnRIoBNwwjYKI31+bKkFQegiadLMFSTKWjDEMBGae+sslEB6ISnPcx54ZGEXlJ1RsCmIYDNUnctHgIDHfCUsNU4AS2EELVKzcuXh/8IYLM0kw59ewEDKeXuEsCGIYDN0koKlwAGDi+g32CVcpu7Vd1VoLMIYLO07JZSru4qgPAK6CJGKdt31wlgwxDAZqku3GcXEmAgKWWDVdCGIYDNUv7nVcsigAHz2AlFK0rDEMBmaZeaxC9wVEF8DtyssA3JNASwWZyRoYA+wgJwFKq2tc0I2DAEsFmSL02Sv8BRHfoq8mzorNqle5tevTg0IYDNImO6KwCizKvvv6rdTA4EcWIcR0EAm6VdqQV1HyOAQ1NuW6S4sk1DAJulubwc1H2MAA5PqdZuS3cR6DAC2Czt9W3dJQDoOGnZbpUANg0BbBZVq9EHCzCOtO1mm2vbNASwWazeYYtnwIB5rFiM27Vp+ImaxU7auksA0HFKCMXt2jj8RM2iRIPxL2Ae5bZbXNumIYDN0lpfoVsdYBwpxNwqZzGYhgA2i9pYqXEaEmAc2V5d5cu1aQhgw2zcLesuAUDntXY3GQGbhgA2TK3p6C4BQMepRnmNADYNAWyYZiAPUgNwJG67WVqlEYdpGC4ZphaLK0U3SsAkSrUa7cqK7jLQaYyADVPeqjEEBgyj3HZthzazxiGADVNa3hYMgAHjbO6wCNo4BLBhGlsl1yJ/AZNIy3Zvr9IK2jgEsGFUZYOVGoBhpCWqVQLYOASwaSp3aUYJmMaybW7W5uFnapp02m2TwIBJlNtu51O6q0DHEcCmsSxODQUMo1RLSr5YG4cANk2jzJkpgGncVo0L2zwEsGmqO21OYwAMI1uVmu4a0HEEsGl2N+vkL2AWKWsVtgGbh1aUpmlWqwQwYBQpRa3KCNg8jIBN025UWawBmEW5pdWS7iLQcQSwadq1ulAkMGAQpdqlxU3dVaDjCGDTVFduN+gFDRhEtRu10jxnMZiHADZNZZVTQwGjKLfVrK2yCMs8BLBp2hulKlPQgEGU67YaZd1VoPMIYOOUU06bBAbMYVnW5kpVdxXoPALYOLuy5ZK/gDmkbW9tNXVXgc4jgI1T2yoremEBBpF2u0mLdwMRwMZpLi2Qv4BR1Po2AWwgAtg4rTvXyF/AIMptbmy0dVeBzqMVpXm2q0q5bAUGDOG2Wq3SSkN3Geg8RsDm2ak0lWIdNGAGJZSqr6/pLgMeIIDNU9kqC+IXMIZlVe5v6C4CHiCAzbO9uCYspqABM0hpyXZlV3cZ8AABbJ7y6pYgfwFTSEvs7LIN2EQEsHncnTVmoAGfeXjRyfZaiV1IJiKADeQ2G6zBAoyhajv04TASAWygdq2hWIYFGEK56xs1AthEBLCBKuu7jIABf3m27EK57dK9klevDp0IYAM1tjfJX8AQynU35zmM0EgEsIGapRLHMQBmUEo1N+5u6y4DXiCADVRZmmMbEmAIabk7K4yAjUQAG6i6sk7+AsbY3Vpv6a4BXiCADVRfLTdZBQ0YQUqxusUaLDMRwCZabyv2IQFGUEJU6vTBMhMBbKKdcpnjkABDNEsVZqDNRACbqLa46LIMGjCAUm5je4c2HGYigE3U3r7nsg4aMIHr7i6tEMBmcnQXAA+45WWX/AXCTylXbS+u6i4D3mAEbKSm22YRFmACS2wubuouAt4ggI1U2dxlGTRgBLe0tqW7BniDADbS1tKiIIEBE9Q2N3d11wBvEMBG2rxzvyVZBw0YYH2jxjZgQxHARtq5c6dG/gLhp9TmOgNgUxHARmrfW9wlf4F9euJpTYC62CilKqtV3VXAI2xDMlOtVdFdAhAa8rl/q5ESqrF0h4vZVIyAzdSsbATpazyAQ1GisrLICNhUBLCZ6mt36B4L7F8gv64qJdTm2mpddx3wCAFsptbGUj1AE2kADkFK6a5vsAvYWASwmVrrq1XyF9i3YF4uUjY3N3kEbCwC2FDrFZdOHEDIKVXdKrML2FgEsKE2y7su+QuEmnLV1v0NLmRjEcCG2tndbuuuAcBRKOW6GzfWdJcBzxDAhmrev9nQXQMQAV6OT5Vw68uswTIXAWyq7ZUGM1dAuKnGzmpZdxHwDAFsqt0tRsDAgR34a6uXy6eVu3F/g13A5iKATbWztBzMjRVAkB34qvFyoklam+u7tNQxFwFsqp2leVd3DUAYBPdZjbR21ulDaTAC2FSl5SX27wP7cLSpIm8nmrY32QVsMALYVI2lxXXdNQA4kvb2CgFsMALYWGvb93kIDISZqm1xEoPJCGBj1baW6IUFhJcSavs+U9AmI4CN1Vy/z3dnIMzaK6u04TAZAWys9urSju4agOAK/vyQrK9ucBGbjAA21/21KhuRgGcJ/hIJd+POGv10TEYAm2tjfYst/EBYKeWuLmxyDZuMADZXeXOpEYJpNgBPoZRqbt/a1F0GvEQAG2zjDk10gJBS7Xp1c4EANhoBbLCtpV3dJQA4pFatsrLIGiyjEcAG25y/p6RiEhp4gcNdJB5fWm5reZX8NRsBbLCdBc5jALzi+Vdbd3mFh0hmI4AN1lxYqDD+BV4okDuSZHNpmTXQZiOATbZ89XpbBvLeAoSet5eWklZ5db3t5VtAOwLYZJWN222GwED4KCFkeXmNZ0hmI4BN5jaqip3AwDOpIyxS9Hh9o2xX7i15+g7QjgA22upChQQGnkkeYR7Z0yloKcX64lrZw3dAABDARluZv88cFhBG7r2FdY4iNBwBbLT1hdtNVmEBYaOEu3Prxw3dZcBjBLDRKku3dunEAYSNbDfWlm7Qh9J0BLDZVu+XjrLMBIAW7er66t2a7irgMQLYbDt3ltttlwQGOsrjb7Wq3dxdu7/u6XsgAAhgs1Xmr7ITGAgZ5bbqi0t13WXAawSw4ea/2dJdAhBYh31A43EXLKHcrWv32MFgPALYcOuVkrBYBw08wyEuDh/mlCx7m5OQIoAANtzu2k2X/AWe7jDXhh/PdKRV2yCAzUcAG669eJXN/MCTlNhbSRXIb6dSypa7WdFdBjxHAJtubXGLVVjAI0opJaTy+kHuUUi5vl5u6K4CniOATbe9OM+RZkCHeX0Sw8q9El+czUcAm27r9nfsZgAekVJKIeQvIXqgoFN7c9fK49Gzu3qdR8ARQACbrr28uKa7BiCIHoTogaLUn2lrVV+b4ySkCCCAjbe9s0w3SiA8lHAra/foQxkBBLDxKgtXWy4JDDzed+MIF4TXg2ClVHP+7n1v3wSBQAAbrz53c4X4BUKkcXeJTUhRQACbb/Hna4pmWIAQUsoHY2ApDrGS2Z+JJClV5e462/ejgAA23+b2PXYUAnsem0A+8FyylOrBJLaXX2iVUisLm8xaRQEBbL72+kpVdw1AEHRqCOvxhFLz/hxHEUYCARwB6wv3+DoNPBjCHu0FpPA4f5WQ20tz7B2MBAI4AjbmfuZgM2BPCJZD3Ftm0ioaCOAI2L7145ZP60eAwFLql/7PR7oYPL+Smsv3Nr1+DwQCARwFd+/f87p1HhB08lF2HvIUwgfz154msJKivrhA+9hoIICjoLx+S3cJgHZH/g4qhR+nAbe3F++wbyEaCOAoaKzfaflzjjgQTI/NPx+SFEJI708xlKK1PH+XRRvRQABHwp25e23yF5Gk1N7mXdmBLpRC+LCIa+f2Usnr90AwEMCRsHTzpwYBjCg6ymNfLdylhXXWQEcEARwJ5Wv/vE8AI5oeHv/7MIKPEsXeX0WqvnJri4s1IgjgaFhfXlQ8BEbEPPmJD8NePLV+96cV3UXAJwRwNJTuzbkkMHBUnl9D6t7CrW2v3wQBQQBHw+7cTbb2I2qeXLjcgfWOdaZgAAAgAElEQVTLnj9KrszdYAAcGQRwRNy9t9AOzzoUoHM6+LH34RFw6dYcS7AigwCOiLX711vMQOMFjPqIKCX2/o3ULycwHP7fTylxxHMc9qe9duuu9++CgCCAI8K9v7ChuwYEnklzJEpKpZQUQkn5MIQf/PsdKkj3zgH2uqVrZf4OByFFBwEcFUt37rV11wAEwiFC1KevJmpp7j4z0NFBAEfFyt0VGrwjGvYGq+LhCiwhpDzy0NXzsa8QQojmwo1NvihHBwEcFbtzP93XXQPgi8dabshHT24f/unhnuT68gRYle9dYw9ShBDAkbF0+3YY+hAAHdXRcavXg2B3ZXFuy+P3QIAQwJFRunOjrLsGwHu/rH7e++2DJVh7f3/4V5XShzXirfvL9/iWHCEEcGTUbt66ydMlmE/+Mu2s9p7bKvXwAa785ZfDvfDRi3sutXlzgSVYUUIAR8f8rZ+bTEIjcjrxmVe+7JF2l6/ebXn/NggMAjg6Kgs3l4za6Ak83a8GvKITj26lL2uwSovXl71/FwQHARwhSwtzzEEjejrxrVP68N1VLd6YpwtHpBDAEbI+N7cVihPZgCN48iMuO/KZl54/Albte1fvNrx9DwQLARwh1Ws//qiYhIbhpBS/GvWqoyen2mtq6SnV3Lnxc8njN0GwEMBRcv/WNbphAYHk1m9e4yCkiCGAo6R67/4GM9Aw2aP9vw/+erCh6zNmq33YBKzc0k83WIIVMQRwpNy98QPPmGC0J4PyYPPPz/inleePbpRw791cZgAcMQRwpCzf/I6HTMABKeF1ACsp6/dvsgQ6agjgSGkvzF91dRcBeEqpDi9YVkJ4PQUthdheJoAjhwCOlpVr32/yFBjm+nX0djCIPV8EvbS0UvH4PRA0BHC0VH+++jMBDPM9+Sk/7KdeKaU6cJrwi9+nsXxvjUszagjgiFm+9XPNpRkHDPbEPmD1YA75MJR6cJaS51dM+/7c7ZrXb4KgIYAjpnbz+nyL/EUEPEjNo41d/bpWqnM37rBDIXII4Ki599O/GnTDgpn2jgJWe+f/Phq3SvHMHb7PJx8msOcz0Pd/vnrH4/dA8BDAUbO5cJPd/jDU3uyzFFLKR4cAP/Y/HdTDJh5e569bnft+sezxmyB4CODIWZxb4BkwTPHwo/yUz3QHWkA/+MXz8a+7c+fHZTYIRg8BHDlbt+6UCWAY4sls/CWQ5REPQVIPT3Hw/nmN67buL9xY9/x9EDgEcOQ0r3/zTZMv2zDLL8PdB6krhThaBEsh5KPX8paqXF/Y8PpNEEAEcPTc//f3Oy5jYETBET/nSnjehFIIIdu3r83ThCOKCODoad+/s+D6tr0C8NZvWm48+oND98/4ZQ11p7taPvXN5Obi3BKTUlFEAEfQ6q3vSv5tcAR8JEUnPtryqb/1zNIcWxOiydZdAPxXsxPDI5LNwDDCE59jKaVU8vGp4wMdCPz4C6mONpN+tuq3f/vXog/vg8BhBBxB7uLa7Tb5C2M92A382N8d4jUeNPXwfqaofeP7b+97/i4IIgI4irYX55eZgQZewJcN86py7efbHNMdTQRwFLXuLFxv6y4COLz9JeMRx69KSh+eAbtL13kCHFU8A46kWiJzLKe7CODQ9heLRzxF0Jc2HGr9X//vTzThiChGwJFUu3b9LkNgQDfltm/9/BMD4KgigKNp/e5a1Y/1JUAoKSH2mmF5/DaqXb3577u73r4LAosAjqbGjX/f9meLIxBGSinvm2Ap1W5szt/a9vZdEFwEcEQt/te/WrprAIJJqb1+Ht5/Q23X787dbXj+NggoAjiiqvcXl5iBBp7Orx4cauvn+S0f3gfBRABH1Z1r/+bJE/A0/j2baV6/vlLz7d0QNARwVC1f/e8l3TUAwaOUEFIp5UcOq7lrt9aYiYouAjiqWgvzP9Z1FwEEjpR7M9B+vFV9fu4aXSgjjACOrPVbP9/huzfwVH70wBLtlfn5OyzBijACOLLq12/e5AxS4BePHyTsyxC4fO32/Kb3b4PAohVldNXyXdNptgIDD0ghHqWw9z0o3dqPf/vPa2Wv3wcBRgBHlyuK/SOO7iqAAPj1nl8lvD8uW7mNjb/9r285BzjSCOAIqyR7JvOHPK0cMMljm37l3hkMnjfBapSu/uf/d4d2OJHGM+AIa1778WqLhtDAI0ooJaT3A2ChGqVr1xfZAxxtBHCUrfx4c9vd59GqgPmUb0+AhWquXJ0ref42CDQCOMrcG1dvcCohIHxcfPXg7dzm4uI62xAijgCOtLUff6wzAAb8ppRamV/c0F0GNGMRVqS5rWzXOF/CgL2Rr5RSKSl9OIfBrX37j2+XPX8bBBs332hb/P6bu7prALT6ZQ5IKaWUP9sCpLgzt0gPjsgjgKOtee3nH1wmoQGfVecX7nIOYeQRwBG3Nnd9TbEVCRH2YMirlHzwix+21u4usAc48ngGHHGuKnSNODTjQMQpIaXyrQm0aP74t29uswMh8gjgqNtNFQe7CWBEmxK/BK8vF8Pyf//Hz+t+vBECjQCOurYoZIdSuqsA9FF7zSf3futH/qrmP/75v+YZAIMAjryKlcmNMwRGdMnHf+tDDyzVWvmvf3xHFyywCAvNH/79fYVVWIgo9cRffXjHdu3u7RssgQYBDCHK1+cWmnSERjTJB78++KsfA2D37jc/LbIEGgQwhBB3rn1bViQwoszHhzCqPvfDHCuwIHgGDCFEs5EbHfJp+wUQREpIofx4ACyUUAv/+o+bZe/fCcFHAEOIitPVW/Tl7gMElj9XgFSt7/71X/c4BwmCAIYQQrjVQmE0TgAjupRP+Sv+d3v3+RVHsuZ5/IksBwgQXkISINNXfWfmjtuz+7fvnt25d7olTGFFSwgkgQDhTVFFUd5kPvuiMJJaBlOkqfp+zmlZuiP6KCt+isiIJ8ROTc3OF11pCn5HAENEci1dQz2unIAE/EVFRNS4VQJL5Hhq/I8NV1qC7xHAEBGpdHYNxwhgNClz/s1t0+rr2fhyzo2m4H8EMEREcpGOB/cIYDQblfO5rzv5ayfnpv7YdqMpBADHkCAiolt7m1xLiKakIupa/uaX3/+x40ZTCAICGCIicrS+vMXGTDSh2t873clfp5RYeveJHVg4xRI0RETEqXR2Pg27dRkq4L3zaa+6UQBLRNSpFl6Pvlp3oy0EAjNg1Oy+W9qyKYeF5mFc3/ev9s7Khz2XG4WPEcCosVc/vMtTkBJNRkXcqwGnpdWPGwcuNYYAYAkap3LSfa/fpbU4wAf0PH/dWYE29vLk/CJvgHGOGTBO6drbpaKtTIHRBM4mvsYY41YJLCOZ5dW1E1faQjAwA8aZktU10BtmCozGpxdHf128haS6ODf7jgkwLhDAOFcMRwd6WBNB4ztLXePqK+DV2ZkFzgDjMwQwzpWks3so6nUvgNt3ttDj3h0MUk2Nz06uVdxpDMFAAONCse3uYC9L0GgStemvSw+85l9NxN/k3WkMAUEA40Kl2Nnx3CKB0fj0dPXZpRIcouWVsdE3aTcaQ3AQwPhMzuoY7Ap73QvgtqkYUdeuYBBxqsdTv73hEgZ8iQDG5/LRlift6tquFMATtdmvurUArY5dfvvyf29yxg9fIoDxuVKlo+uh5dq+FMALp0Ho4hHg6vrYzELZlbYQIAQwvpCL9nT3ul8kF3BPLX/dXIE2xXicBWj8Cac+8YXKu+l5/qKOxvFFbTf97GfGrUuARYwkEhtcwoA/YQaML+VjnQP97MNCo/hiNedibUddKwEtIk4pPju76VJjCBACGF+ptkcedbIEjUZmRNTFFy2VTxPxJWpQ4k8IYHwlX7pz9wkvgdFgLvb2n9+A5FYJDic7NTG9705jCBQCGF/LhXsG2ynHgcby+eLzaQFKd55xdSqrY9Pvq640hmAhgPE1u9TZORJhDoxGpPLFXUguNKhOav4fi0euNIaAIYDxJzkn0nk/wllgNChjjHs1oI2U52bG1213WkOwEMD4s6xpa31EAKORufZ4O5+mZl+fuNUaAoXzJviz/FJH67+3et0LoP6Mqnuvf0VEpLi8/IEFaHwTM2B8Qz7cN9wdVubAaBx69p27+Vt+Ozm1xC2E+CYCGN9S6eq5305JaDSO8/x1NYDV2Zsce73rVnMIGAIY31IqWeH+OyQwGoOeF8Eyrt0BLCKidn5i/Ld1bkHCtxHA+KYTp/XOCNcioYHUnmXXbkASUdXC8u/j7ysutYfAIYDxTZppufuszcXBCqg/FXM+/dWzYljuPdKOfTTx9z/YAY3vIYDxbZVq653BmGunJYFbcPr41nK3lsAurj+L5F5Ozm641R6ChwDGd2RNW9uDEAGM4Dt/iN1d0jH2wmT8Pbd74rsIYHyHZsJ65yEXRiPAzm5gMKe7ny1X81fzMzOTHAHG9xHA+J5yMRYZvsMMGMFljBqprT4bUZcnwFJemphbpgYlvo8AxndltK37UcTrXgA3YmobsWrvgV3MX9W9mfG3TIDxAwQwvi8f63vYxRQYAXd29YKLB4BF1Cm/nRhfddxrEcFDAOP7KqWOjmGOIiHATC11azcAuzr/raxMxBez7rWIACKA8QNZp727N2wRwAg0dbkApYiIsxePz2272SKChwDGj5xIqGfAcnnoAupEa/ufVVxefxaR/ZmpueWqq00icAhg/Ei10NLzqI38RTDVQlcvfugSdcpzM/F31MDCjxHA+KGcdPU/In8RXKfbr1zNX60cxMenEy42iUAigPFjufbYcCvlOBA8p/dZqxqX3/+qVg9GX7zadLFJBBMBjB+rVKLmYRtzYASQUTEe7L8SJz03OvOBEhz4GQIYP3Fit7Y/piQ0gkRrZ3+1dhGvywfpVAuzk6MfOIGEnyKA8ROaMV1dPa4W0QVu5uwvjKa2+uxu/kpxdXL6zaGbbSKgCGD8TDXX2TUcphwHgkblogqWe41qdWs2/mrdzTYRVAQwfqpQCVkPo6xCw6/0W8+mqhEVdX3+66SmXsQ/cgIYl0AA4+cyTqzjIYvQ8KtvP5mnNyG5+9iaajY+MbZccLVRBBUBjJ+zM5H2oXYSGEGgp5f/GjHq8vlfEdX8+3+MLuRcbRSBRQDjEkrFqPVrhPxFANQOHRkVD84fiVNeGfttKeVuowgsAhiXcaIt9/rCXvcCuCxTezHscv7apeTE+PyWu40iuAhgXEou1tbX53UngJ+p1X0++8bl/NVqdvJlfI07gHFJBDAupZKPmGcRSlLC587e+nox/1XJvRqdeld0t1UEGAGMy8lVWtvuRziLBH9TI7VCWO6//1WtLsZHl5LutoogI4BxSRmJ3usOkcDwLz0tQile7L9SUz0eHZ3ac7dVBBoBjEuysxrq7Hb7WAdweea06oZx+/4jERFxjsdfzq2r280iwAhgXFbpONLxNBziNDB8SM8nvqfcfkxVi/MvJ96VXG4WgUYA49IKpbA12MoUGD5kaqvPerYL2vX8leq7id8X0y43i2AjgHF5aael6z6vgeFXRmuVJ92/OUS1vD0+ObfrcrMIOAIYl6fZaHdPFyUp4UdqzGkJSrfrP4uoOofx8dmPvADGlRDAuIJyLhwaauc0MHxHT9edVVyv/yyiTrXwemz8PS+AcTUEMK4iW411DkW87gXwZ7X6G96sP9vF7YkXb09cbheBRwDjSjKh6L37XncC+JKKMWpE9fwkkrvNV7IvfptMuN4ugo4AxpXYhc6WRy0sQsNP1NT2P3sy/xVx7Pyr+KtVXgDjqghgXE1e26Jdd9iGBV85fyA92KOvWn0/FX+Xdb1hBB4BjCtK2yJ97V73AjijclGHw4szckaPJ6dnt91vGIFHAOOK7OOqFRvmLBL8obbwe1YHy5Onsvh6fHql6kXLCDgCGFdVOQ7H2vsoSQmvqbm4/1eN8eD8kYiI2B/j8TfsgMY1EMC4snLaCvd1eTXdAE6d56/W7kDy5nnUrYnJPzbZgYVrIIBxdYWMaent4GIk+Icnx49ERJzs+OzEStmTthF0BDCuIZsKxZ6GCWB4zchp8Suv5r+SW4xPvsp70zaCjgDGdWQrYbuPw0jwlorUDgF7cvxIRETzc1Oji5TgwPUQwLiWlG1FH0RIYHjPnH/jOq2+mY6/3uAFMK6HAMa1OMfRijUSIoHhPjXnly/o6e1HHj2IevD76Mstx5vGEXwEMK6nkg6FWgYtEhiuMxffezj7FRHdefH7q0/kL66LAMY1FfJR7exnIxa85tkj6OQmX4x/ZAM0ro0AxnVl0xF7sJN7GeA2NbVNV16e/hVVKc+9+G2ZDdC4PgIY15YphM1IlDkwXFY7e3T6I68eP9Xqymh84dij5tEQCGBcX6oSjgzGKIgFl+hnz5oa8fD0r6g4e3O//bHpUfNoDAQwbuDoxJGnFjUp4Y7T1Rat3f7r4fqzqNH8xMTYmu1R+2gMBDBu4igTjvWzCg03nd2/4OH8V8TkFsbjS7wAxo2Eve4Agu29JZ3/I8IUGO64KHnh7bqLke13f7zjCiTcDDNg3EyyYDtDrELjFqk5//6zxRZPnzjdmYxzAhg3RQDjZvQoq529EVahcXvM59+f7cTy8olzMjOzYysFD3uAhkAA44aco3w29ozjwLg15/l7ugBtjPH4Lsz067mpmYyXPUBDIIBxU85xONoxQALj9uhnZ389u/nonBbm5yYX9rztBBoBAYwbq+Zj1oNO1qBxW2pnjs7z1+sNB/bi9PTcOi+AcWMEMG4uX24J32v3uhdoWMacrz77IH+dg/hkfK3ibSfQEAhg1MGJ3RId5m5C3B5zdgGh19ufRXbiL2dWuIIBdUAAow70ONLW0R0hgVF3amor0LVrf9Xj3Veqmpl8+fv7opedQMMggFEPdqpSivWHvN4dg4aiRlTM+Z1HxvvVZxGTmh6deJfzuhtoDAQw6qKUrLa19lskMOros9Q1Ih4vPouIqGQWpicXUl73Aw2CAEZ9FFNWrL/T8n6MRMM4e+er4oOXvyIiKqXFV5Ovt7zuBxoFAYw6KWYcaevztEA+GoOaL39yWvnKBw9WdXlmdoYDSKgXAhj1kklrW18Hc2Dc2Pmtg2dHgC9+0VPOp5mZufdsgEa9EMCom0zelsetPhgnEVjnZ41ETotfqX/yVz+9mouzAQv1QwCjfk5CsVAXBTlwfefrzFqrfXW6/uzx4aMae3dicmz52OtuoIEQwKgfLRqJPAr7YKxEwGmt9IYPLj46p4k3Y+OvuIEBdUQAo46K+aiRh2Gvu4HAOy0+qWr8MfsVcTLxsRdLWa+7gYZCAKOechVjxwZIYNzc2clfX8SvOOnZ+Oi7I6+7gcZCAKOujotWKTrkk0ETQaSfbcLy+t7fC7nFiZfTSa97gQZDAKO+jnMhK9bNxQy4LnN+9a/6JX3FKcRHXy7te90NNBoCGHWWLptQ+112YuHGfFD6WURExc7+ER9/s60//1rgKghg1FsyU03aIxTkwPWp+Gf5WdXJvfnHyz92KICFeiOAUXfHmZCEB8IkMK7hdPHZL5uvRB07Ozn+4sMu+Yu6I4BRf+mypa39lk9GUASEXhTh8M/uZ1X7ZGF0bH6H9WfUHwGMW5DKhpzwoOV1NxAopnb/rzFi/LL8LCqSm30xusj+K9wGAhi3IV0wTqSfpwtXoCLGnB//9QVVLcxOjH/Y9rojaEwMkbgVqYLkIwOcRsJlqYiIEaP+uHhQRERUNPf+ZXye97+4HQQwbkcyo9niYMzrbsDn1Jz+c/FLfolfUSPFV+MTi5vkL24HAYxbks6Winov6qPxFP5Tu35QjR/zV0RLC5PxhY2q1/1AoyKAcVtO0k7Beuaf9UTcJhWjV83O88t/jRojxlelJ0VETPrt6MT8etnrfqBhEcC4NfnDQqXU3uGbEyW4RacJep1/5/TQ7zX+A7fKqSTjY2OLm+Qvbg0BjNtTTuSKcrfDV7Ma+I9R/5z7PaNaPnodj78lf3GLCGDcIns/VS7e7aYkR5PTbz8An61Z+y2A1anuz/z3y9fsf8ZtIoBxq1K58nH1XsRXgyvc9s0/fhVzvvfKd/krxZWJ8fjHhNcdQWMjgHG7Usl0of0+B4IbWe0Y0ZV3YH32b/jt8dDqu/jozNu01/1AgyOAccuy2ZboQCer0A3MqJFvhOh3Fp5Pf6tW8coY8VHhjXOlpanZmZW8191AoyOAcdvyOTF3en1ytytuwXcuT/jBH7i5+Mdvq88iIuW18ZmZ1azX3UDDI4Bx6zLJYutwjL3Qjer0Re6P/ni/u0Bt/Dj/1cP5sanFgtfdQOMjgHH7cieVfKUn5ruBFnVkfrDifB6yZ1+jX/6yv1TWf385sUL+4vYRwHBB9qRYtAejvhxuUReXXUk2clH32Z/PQ2lpKj71Pud1N9AMCGC44eS4Ih09Ua+7gdtSe6F7PglW+TJeT5egtXbwSMX48tVvzev45NQS+6/gBgIYrsjlxKn2sQrdiL5YVq795OuazsZ89vtqTK36sw9p7s3o9OxH8heuIIDhjmyuWpWuFsvrfqD+Luo5/2Ba+9lWLd/Of51KamZq8hXvf+GSsNcdQLPYsU207T87ve4GbsHFBqzvxKqKnO7Acox/81dKhxNTE58OuH4QLmEGDLfkMsViuStkMQluPJ+d6/3xl/nw2oUzWjlZ+X10cumI8s9wCwEM12QT2ap2x8J+HYFxfeaL777/Bafrz35Uyay9+H+TlL+CiwhguKe0nzwqxXqVmhyNx5ivN159+bt6+iWWX//sNfn6v17Ob1e87geaCQEMFzmJdDnc0x7y7SwIt8y3f+6OvfTy5dImy89wEwEMV50c5ctdvYYEbja1Sxd8+6euTuHl/3m9qz//SqB+CGC4K1ex7NBDLkdqOj5OXxHV3PzfZ7Zsr/uBJsMxJLhsI+aUWv854uPRGM2nuDT7fpfjR3AZAQyXOcvhqDj/QQDDRz4uLmyceN0JNB2WoOE2TWVyWacnxLMHP1Ax+Tfx2dk1NkDDbQyCcJ2TSpcLTl+EnVjwnqqTfzcxPfeeA8BwHQEMD+T2jkp2TzRMAsNbKiLJyYmpV2vcPwj3EcDwQiWVKZdaO0hgeEzt1Yn4zNtN8hceIIDhCSeRzJlov6/PpqDBqYhU16Ymx99ulr3uC5oSAQyPpI9LhXJHh/i4OhIamoqYk4XR0fhK0uuuoEkRwPBKNl2qlNu62IoFj2h5d3o6Pv8x63VH0KwIYHgml65mCoOd5C88YYpv56bGJ1l+hmcIYHincOw4+fZupsDwgJN7NTk28+GA+s/wDAEMDxUzpUq+o5PK0HCZqp15PTk1s3LsdU/QzAhgeKl0mLYrfR0hEhhuUqean/ntH3MbLD/DSwQwPOUcZwtlq9diKxbcoiJaTcTHX77fYfkZniKA4S09ThSkrTtkkcBwi1Y/ToyPvzryuh9odgQwvJY/yhWlq1U4EAxXGFNenJqLf+D1L7xGAMNzxXROylZ7hACGC1Qy8xNzsx9SXncEIIDhveJh/uhAelq97geagDrHs9Nzs0sUf4b3CGD4QDWVl7LejzAFxu1Sx157MTo+/6nkdU8AAhj+UDkulUuhnih3M+AWqdql5fHRmffbttddAYQAhk84R+lCuTrQYnndETQsFa2UVsZGf/vI9iv4AwEMn8imj3O5WLtl2A2N26BqnNTs+NjrdZaf4RMEMPyimMiWIqHOsEUCo/5UtLofn5x89anidVeAUwQwfMNOHGWPT7rvCgmMujNSXZiYis/vOF73BDhDAMNHMplsoWB3h3kTjHqz8/Mv4nPLCa/7AVwggOEnmWQ+kbvbS11K1JWKU1yYGJteznjdE+AzBDB8pXyQLRWKd1uZA6NeVMSu5Ef//l8Lm1Wv+wJ8jgCGv2j6JJPP6Z0Q9yOhLtRRp3w49XLizT6XH8FfCGD4TW5rP5Gu3m1hHRp1oGpr7uPY+O8Laa+7AnyFAIbvaOookTg8iXWqksG4ERWR8urs9PTUGq9/4TsEMHyosJ9I5EqhOxFKU+ImVMTJLUzMzr9Z4fIF+A8BDD/Sk+3DvX0djBHAuAFjTOaPV/OTb7bZfgUfIoDhT07yJKvVXopD4ybKu6MT8derabZfwY8IYPhV7sSpalsHq9C4JtXc+4npmbmNotc9Ab6JAIZvlY4ypZJ1N+p1PxBIKnZi8uU/JpeSTH/hUwQw/KucyuQyhXCrYRaMq1FRza9Mj8UXNgte9wX4HgIYPlY9PEqliiGqcuBqVFWP/piZefHm0Pa6L8B3EcDwtezBwf7eid1hKMuBS1IRI7kP8zOT0+sc/oWfEcDwt2rq4CBTlvaoxTo0LsWIOIdv5uanF9dZfoavEcDwu3Ji6yAd7my3hHuCcRnGWZlfjI+9OeTqX/gbAQz/K6Yz5VK4N8wcGJegmcWp6fHFDaa/8DsCGAFQTuYKTrifAMZPOdXk/Nzc3Juditc9AX6GAEYQOMlMNW/3tJDA+AE1IpXDibH/O7uc9bovwM8RwAgEPT7JHqXtuyFKU+K7jFZTs2MvZ5Z2OXyEICCAERAnh+lsttwWM2zFwreoUS3vzU7+PvXhxOu+AJdCACMoyocHiWS62BIOEcH4mooRe29m/O/jb3d5+4uAIIARGJo9SiZTqVJbyCKC8SWjTm45PhWfX0tR+hlBQQAjQCpHn9a3nFB3xKI2Jb5kFxZmXo7N7ZW97ghwaQQwAsU+SSYPDgt32tmMhc9oeXfstxd/bLD5GUFCACNgSvuJo7xtdYa97gh8Q+3S+uSLicXtktc9Aa6CAEbQ6EkyX8qFH7AGjVNaXHnxj99Xjnn7i2AhgBE8pVSqkC+HYyEyuNmpiDrlvcnRsQVKTyJwCGAEUCVxUizliu0hilM2NxXVavr99PjYwhbLzwgcAhiBdLKzvnd4UumMGuVIUtNSVSlvTY3+9+z7w6rXnQGujABGMFVSB4eJdFrbwsKRpCalos7RwtTE9NIWu58RRAQwgqp0uHl4XK7/Im0AAAymSURBVNTu2i2FZHCzURGncjA5Pj63mGD6i0AigBFc5f2Dg4ODbFuH4V1wk1EjIk7y9fjLyYVtdl8hoAhgBFn2MJnMZk0bu7Gai4qok1udm574Y/WAm48QVAQwAq16tJ3KFyutLZZRlqGbhYpK+Whhdmw0vpX3ujPAtTFkIejM/YfPf/nlX/8SDQnz4CagIupUttY/Ln3Y2Et63RvgBpgBI/CyO9u7mbJ2hLinsAmoqlNOvpmfnZxf2mb6i0AjgNEACvs7h0fpaneUKXCDU1FH8ysz4y8n/9jJUXoSwUYAoyEUjhLJ4+N8R4wEblwqourk3s+MT0yvbmUdr/sD3BABjMZQOTpIpHLFLibBDUtF1akkX02NT7xeSXH0F8FHAKNRFA/205njUkcLCdyIVESluPtmamJibu2I2S8aAQGMhqG541QidZSJtTILbjgq4lS33sxOTb9Z5dpfNAgGKjSU2JNf/+k//9fDMBHcSFRExDnefPNuaWUjw+wXjYIZMBqKnTg4SCZOrM7a3y2J4QagIqrl9NupiZezH7azbH1GwyCA0WCKB6lk6jhbtKKGa5IagYrY5fT7+amZuXfrR+y9QgNhgELjMb1P/unJ8ONfH3rdEdycisjJp/dLS+93jypedwaoKwIYjSjSN/T46a//8Txm8YgHl4qoarW0+e7D0tpOIuN1f4A6YwkajcjJ7qYyhVwxEuOmwsBSFbXLhfVXM1NTb1YPyl73B6g3Bic0qlD/yN/+9i//3h0WEZ70wFFRdaqF9Q+rH5b2jgpsfUYDYlhC42p98MvzX5//rSfCbqyAUVFHnOrRxtby+629vTQ7n9GQGJfQyGL3n/3T/3z6tC9qed0TXIGKOraTW//wYfXjerJE/KJBEcBobC33nz7/5Ze/PbZ41INCRcU4ibWN5cWVg+SJ190Bbg2jEhpd24ORx3/92z/3xEKGBz4AVMSpZlZXP35c29mn7BUaGeMRGp91/y//8h9/fX43bAwZ7G8qIqLZzdXlxbefEpz7RWNjMEIzaLv3+Nlffnn6PMa5O/9SMaIqdmZ9eXl5bfcozewXDY7xCM2gcrx7eJg6KTrtvAv2KxUR41SLH+fnpmcWPu4V2XuFRsdohGZh3X/y1+e//tu9Nq87gm9SNeKktzffLS5uHpZJXzQBAhjNo+3+8OO/PH76L3c4lOQzKiKqpZ2tzY3VTzsHSeIXTYEARjNpuT/89Jd//+d7kRBXJfmIijp2+WB9bW1jff2o4HV3AJcwBqG5hHsf/u35k18ft1uWJcInwHO1fc92dmN1bWl1O32S97pDgGsYftBswg8ePXr+dOTBYLvFB8BrKiqq5cSnjdX19d2DY9vrDgEuYvxBE7oz8vjZk6e/DrVyVZKXatcNOuXUp7XlDx92khz7RZNh/EFT6uwfefLL0PCz3phI7QQq3KUiKmKX01s7m6sfdg+SvPpF02HcQZO6c//R4OCzhwNPuiIW9bE8oKJ2aXtjY2trd3vnmNt+0YQYdtC8ol1PRkb+9fmzrtN6NHwa3HG24FDe//Du3YdP28Wqxx0CvMGQg2YW7ep9+nhk6MH9wQ6vu9JEVESkmt7eWF9a3Uqmil73B/AIAYwm197/aOjRowcjD/rCbMlyg4o4duHgcHdjdXV1n4LPaGKMOGh6Vnvfk+GRZ0+HBymNfvtUpZrc3tleW149ShWIXzQzAhgQae+59+jBvafDjztaQxaFKm+TU0qsrn3a2D44ShSoOInmRgADIiLS0vdoZHjkybOBlpgxIspHo97UiOOc7O3vLL9b2U2w7RlglAFOmY67/c9++XXkSX8rn4s6Ov+7jJM/3t7c+Li8u59h4xVAAANf6Hv4ZPjh8NCz7ggL0fVlV/d393a3Nnf29o45dgSIEMDAV8zdoefP/zL0uL/d4uNxUyoiRlTtQv74aPvT6tLmXpF9V8ApRhjga119j4YfPxr55V7UMsbwOvh61Kg6IpYpHx/s7u3u7R8k06kTblsAzjG0AH8W6bs/9PjpyMjD1mjYEj4nV6cqoo46Wjna2tnZ3No7TKSr7HoGPsfAAnyTdff+8+fPHj8ebAudlU7k03JJKqKOI2prJr21/v7d2uFJmakv8DWGFOB7uvsHHg0PPxwauhvzuivBoSLqiIqIndlf29re2j44OmLTM/ANBDDwAx33RkZGRvrvPWmNWFSq/Bk1taVnW+1K5jCRSCwvbx4cc80v8G0MKcAPhTp6h4eGnz1+0tkW5ePyIyoqxhGxxEnv7Xz8+GE3kc5VWHoGvocRBfiZaE//w8GB7t6BRw9bYxEmwt9Q23KlRlSLh4nE7tb29t7Bcd7rbgG+xlgCXIbVem/o2bNfHj/qjISN4YPzJRVVrTqO46QPkjtbK2ubh9yzAPwM4whwSVbXwMPhx4+HhgeiIev0s8MHSEVPv7Uzn/b3Nzd2k8fpTNbrbgEBwPgBXF64b3Bo+NHwwND9lrARPj9ymr6OXUrtJQ42d3d3DxMFKk0Cl8IAAlxN6+Dzx4+H7o88bvrbg2t1NYxqqZjc3vn0bmUzSfgCl0cAA1fV2t0/+HDo2bOnd2NN+QFSIyJ6OnpUMwd7W3vbe4fJZOqEUlfAFTTl+AHcVOz+0MOhob7uew/uREKhZtoYrefHfY1Ru3iwt723ubGzl8qWvO4ZEDRNNHAAdWVaex+OjPzl8WDf3WiT3F14ut3KsdRWsUqVTDL18f3S1n6mQrEN4OoIYOD6uvoeDPb03bvXP9DTGfsqhRvoEqWvVpZVK9mdvWTyKJ3J7CcOk8x9gWtpnDEC8EbrwKPhwf6+rtaO7oE7Icu6KFnZIJ8uVRFHjBijIupUTtLHmeT29vbOfjJXotAVcG0NMkQAXoq2tHb39A7cv9fX1dvb2RE2qpbRs4PCgf2QqYhRFXFUbbEsU7ErJ+XS3s7Wp62DTK5QKFJrA7iJwI4NgM+0d3Z1dXX1dHcPDAz234nWdmZpIANYL37gqBjRaimzd3ScyhfyWk0dHh4eZThuBNxY8MYGwM/Cd/qHhx+MPLrT3tHS0W6sQFatdE5P+Irati2Vykk6ubO1vrGTypYcx2HeC9RHAAcHwN/CHe0dXR3d/T09vQ+GOu+0XhxSUnMxufTVR++sV1r7gTq2o6FQqFwupI929hN7++lMJneSY9oL1JOvRgGgYYTu9nR3dw/0xDr7enp62sNRy4QsS1RVjBEj6vXZ4S92NjtiTO2vByoijl0t5LcOM6FCvlTI7u0dHR4V2WwF1B0BDNweE+noe/Do4f3Ou/cidnt7ZzgcVrGMdRbA5nxS7PYnsTbXVSOiamnFWKFaf+xyxSnms5ubW6uf9o8LtrLkDNwWAhi4XbHOzs6Wljshjbbf7bzb297W2dPf1mL98LNXzzPEelY1UkUu0t6pldRQNcayjIpUy7liqZJJHiQSJ/lCJn2SPuZKI+BWEcCAW8IdvX39nR3tvd2tbR33B9pClrEsYz57R3y2+emSp5e+WEb+3terqBrz+dZmY0RV1VHHtm0nWzgp2uVypVgqV53jw53drVTZVqo6A7eOAAZcFQpH2tq7+u89GOzraG1p6w6FTDhiWZYVtk53GBsTsr7xhth8VZCq9sb2PFmNfP+t8pcTajVSqTrlarlcyVeKeweJnYN0JleqVB1H7FKlXI//SwA/RwADHoh1dHV1tMaiLa0mZLXc6eiItbS2Wm2dLaGQZUXDofC3L3g4i2Bz/nNzcS/Rd6fAtl111BgVEbtcKmTtcjadTmXyFbtil9PHJ+mTXIUXvYDrCGDAWybUdre7q+POnTvhls7WWNSyWqPa0xmNxmLhcEhCcrpX62wOXFtQtkJfV2iu/cdOQ1pFnWql6FQrjp3PFbJlCYeqVqhUKlVKxUrp+PBgO5Gvba9isRnwCAEM+IGJRCMmEo2EQsaKtkS7ujra2mLRWDgcCplwKGxCIYm0hEUsY6ullfJAt6VVYxyp7bJyjBFRY1nqOOWqcUr5TLqYSRULxUIhm88Vq07IqBHbVse21S6Xil7/DwMggAH/ibbeudMSi0QjoXDImLBlWcYYK2LUGHXEaLXc3WmcihFVMaKOOlpbirYcdcqOpXa5WCgVcqVSuVAsM8cFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAgO/5//dklgqEntRTAAAAAElFTkSuQmCC" height="1080" preserveAspectRatio="xMidYMid meet"/></g></g></mask></defs><g mask="url(#bac4022113)"><g transform="matrix(0.75, 0, 0, 0.75, 0.00000622222, 0.00002)"><image x="0" y="0" width="1920" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAB4AAAAQ4CAIAAABnsVYUAAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOzdy49u2Xke9ue9rLX3V3W6mxTVpCRLCiLRhmQidgAzcRQksDRIAgRxggzEkR3AyEBA/oLMQv8FGcd/AjP3wEhCJgigRGlObEp21LJupiirD8m+nKrv23ut95LB+k4rMXKXxCap9wd0N5o8dU7VrjqNOs/34HmBUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFJKKaWUUkoppZRSSimllFK+f9An/Q6UUkoppZTyyctM4GvAy/fee/ny5dv45ptvnyeAl9uGn/zo7bdffvY833v59suXbwN4++2Xn337JX7qIwBEX379tm8DAL7wL/zMRP+X33Jn5re+/vVvPz2993u/9/7l8qUvfenP6KMrpZRSSinlk1IBdCmllFJK+QH2zjvvqJ6AMU5yJwskMiJBiUQmIhFBADMJCxElQETMJKzMTERE2F+89dnP/zXg7wL42tf+BoBffPkSwNfefhvAL/7ifw8A//Vfvv/ry5f45d8A8O13/6I9vdnf+MyPfP4XgL8L/Bf/wrv3z//RV88PX0bEmNPDgQTII6Z5Ih9+5Md+/hf+w6//vb/325/+9Kfl/c623m1hZhEmYmZhMAuTAOpCHw0eiY8+QqXVpZRSSinlB0IF0KWUUkop5fvOO+/8VxEPcKV4ECiLCMCZQsnEwsxErMQCR/v2+bjvr9wHT+dETgdJpIE4EhyWTpnWVYiViTMjKBs1acRQMBGlAJEOSgFnJBDEgkx34yQSVqYIC4DIiRiZ01wpuTdYZobZbK1RpgMxzc0CQcGkHOZzzttxtk2E+Dxtpru7qBzTr+dNWUhEWad7AqqsLGAl8sbCAtDWks7U8YhvfhM/+xnfxMf06eEREemRkQgAEJAGKzSS0dr8pV/6O5/057OUUkoppfz5VQF0KaWUUkr5JOVXvvLd3s+OVy8kNJMoI4PPs33X/W06uPWNmQH0CADakr1rQ1D0pswgEJh1a0i4JzMRgEjKzMwkj+mB7KyiLKzmHh68cuWmrAIPNyM3IlLVCENGgigzIpiIQEgEnDxCQoiJ4DaJCcwMApDpSKIkMDLS5gx3Zm6q5uHTxjhbbyIameYWibb1Me16exZRYlYlczhSiJmASPdgAot6WlgACOJMWOacfsyYNpMoLMwRlBEJVsqWyie1y+VZxwZnDrkZ3v7xn5bHxy984f8wEvJ/sxBSSimllFLKn1x9u1lKKaWUUv5sZX75/W+9fT7vr77zqQjKNYcBJoCSHs74C++dv/Xihb85aed5SxFJmu6RREzorXdtRBCCMpqqqAqJKksTRXpEpvO2MUB2JggJuAGRERmWmUiHJxGxKBEifJwnQCyq+55ucd7CjJm0dWQi3N0zMwElzkx3zwwgQEGchEwgIjJTWUSEhMc5wl1EIiI8bBqTqIp7ZCYBkcHM+74nEIC0BkKGZ6ywHNIbqyCBCERGJlhY25wWkQAnOJiD+Hba0/VIokwious5bMwxHCzEMpEJEm4kLRzT7A288du32y//8i//43f+h8j8wr/2NwD8w1/771599yUREUIRn/nOR4+38blvvk9f/vIn/VVTSimllFJ+SFQAXUoppZRS/nR89atffVNnI1xkEgVTMEEYl7eePvP5d3/76385zmZIMAFgUUoKd2VhYSY0JhISShaoqBBxIsK1KTHnnDGn2WhKDGRkkhMgyuHT3aSpMjPBpoVbuBMRE4kwQMjMiMwEUrURUYRHRCaYJdPTI8yQSUQiAsDmzNcF4fBwt8wApXBGeGYwk4iwyIqhVx6NTIAykJ5EAIhAHg6AiUEgAhEnMtf/ue4f3v9KEBMTEsjXmInFIyMJxJYIsLQepOEEJhAz8TRzC4B779I6REg0IcPmeYxjWkAB8QgkBTDCI4IZlFCiYBIbF4m/8qu//e7Pf+6jNy8BWok9KJXx6c/91OPjpz73s3+1GtOllFJKKeX/k/r2sZRSSiml/Il86513Rh4Gf7bx3UN/8nIjF7QbE7GRdohkYsXOZI4EhFtvjYTDUoiYw91BqZIxJ2MqsxKE1vgFITPNfJ42h6ggI2y+7iMnkEAyrzAXyBUmGxJrUmNFuuEe7hnJKkSEzI/z3/AID2GmREQQ0T14JopMs4kEMRMSlEC4W0YQiPUeQAMgJndfiTaSkchMImZicyOQqkQmEswcCI/MDCIw8wqc1y/9xwlvIgkgSuIAJSgTHhlA2zaCRBKJZMLD0gOAsAqrNCVpYEmweVpSJFR2iM6IAGXycR4ZqSqJpHBkmJ8YbunJzBEDHMSwlNZSxu70V/7dv/0b/8t/2979p5fr+ZN/8N1qSZdSSimllP83KoAupZRSSin/zzLzvd/93fP86Onbf0hilEzCjUWaKHWa+1N+YEDGyemc0VU2SpV88bDtvYEjzGOOzJhjjjG21pjII93DYppNEVIVsymUW29wZ+K+7WkOM2KiDERAKMP9PIky3I7j1rr23jx8jHGOue8XIj7HaWaZKSLMnJk+prtHpGdEBoDeuqqa2Zxm5i8eXqjonHPOSUSPj49JmGbPz88i8vj4KCKZOed094yMjMwMJDOrtm3rt/OMzK3vzJpJ5zFFtPc+5yCibdvGmJm575tHTJ8RzsytrUZ2mJmIiMjr9JtAnESRRCwJsnAgidFai4jptm17RFyvVyQYWA8pM5MoExEZARCJCiAETuIEIjOSRKT35uZM1HqP9Ok2jhFJnnwAY+YMp9QUJQIxJUDT/vqv/dY//kuf++DF7rHidGYmZgD4N/79v/XJfqGWUkoppZTvNxVAl1JKKaWU/3Pf+MZXer7gpB798vjmj37+i7/+ta/h8bpNmuISvW3ShCB9a6oKcLBNzDPnaF2ZMuwMmwzbeidYuhEo3OecqsoiIE5kZPicQIJgPgkpRIjMiHDAIyMog4B1mc9sjvNgIhESZSLKjDFHAsJyuTwS83GcEQ5AVUGUERnBqn2/nLdruIlo651F0j0SCVZpTBQekQmCimSmZwQRMSsRMycoiHzONEMCqtQUZkwkKhYBEGsjkgyM2wlAVGkdRsyMSCJqvSfgGWmThKV3MGdEmqV7RjDzvQpNDFaIYu1QzwEECESUuM+JRMQYQ4SJmDzWmIdHgIVFYxoAVr1/35/I9U9mug+McGaGOZhAcEckOVjaNpOmGbixCiCJHLfz1fPTHJbM54hEAprg3gGgCQBEkiUliPoUNX6cX/zir3wSX7+llFJKKeX7QgXQpZRSSikFADLz29/+A7s+PX3wnpiBAjyv+uqN+PHM6xaScPNMIk8oo2tT1W1r0pVFYhjsJvaU4xrzpqqEdJvnecvwh30nAjKY+OOqLwmD5b59HOlrudkNmSsIdnMbxljtZyeAiTPDbI5xStPe27ZvGT7nnG4s0vu2bTuBxnkmEZiVGZmZAZD2vj08nM/PYdZ6Z1FmynAiAQsSGZEe951mooiIDKgCoHAQE3MSp3uaEzJVwZLjBMDCK1K3TCJGUoyRa7xDBEQUjiQwkQjWWkgYMVNrjsxIcg+zDL+vRYOIBSxBwiKU6TbCbb1XzKzKmYgId2dmAjJCmJl4zkEs2reYE5nSWmaGe7oTE4vE/bEHawvP2/V57VlnwgORaNseSeeYEGVp2jrLDqbnp9tpFqDTwywdsUZVOEHCZhkRyXq4dAz97LO92jn6dZIFf/cJX/rSlz7hL/RSSimllPK9VQF0KaWUUsqfR++++/fz0EyFK4mq0OMbn/rsT/3cP/knv3a5HsYuEUzoQr1zF2pCjZDpyZxMeYz0mZFAZriZpQ+EbZoUFj6QASSACCdQb32d1QPgZnNMUQXBI8YcEblfLtP9OE9zJ+be2zzHCrz3vm2teTiBhFlFQQj3/rDrvpFIzJlzUlNSJZX7UvI0XC5ojcaA+1qhJhABOQ1I9E4Z8LiPQRPD3W3O8wTALK13IN3sOI6IFGYWIULEmvWgiPuciNlkQu+97zsIz8/PzKyqqgJCRIw5mflh22PJXP8QFiIGcJzHCpFFRIQBrIkPZonIOaxvXVWQebvdjvMA0HvrvR/HaWZA2rTV1X64XPZtvx03gLR1m0ZEvW9mc84x59CmfWtjznU7cWstIp+fnrS11loEIuCJ+96IO7OyiLAwKzEfw0CkfdsfX0jr5smtsTZVSeAw/+Dp+RjhxB5IYgKDqXf9rX+OH38LyumRhJRu3Iz3Uf3oUkoppZQfbhVAl1JKKaX8uZBf+cqrT3/aN7m+eQl1EzO9xoeXkF3bFGzaqCs1ZmYgJrkhfOtKmTGPGFcahzJoDTWcExnM7G5u5uagICSTEwUQiFiLE0xMzELs4eHBzAAyk5gABNLdAWrbHpnmniAW1iY2ZkSyqrauIuG+GsEMImRGSFMwmVu4U0B7IxEQuc1wp8hUTSI7T85kWhcCk0DKTExBBI97KTvTw1e6bHMCIGZtysTIPI4jItY6MwB3XwMZibXQEYlkIhEmkcw4xxAmUSbme6naHUhhiQiPCA93zwiVpqoicr1dzYyZmYVA5oZMEJg5IuawbeuqCmDMYWYiuratz+OMzNba2hjJzNaaiMxpwtK37TzOyGitr6fmbqKiKnPOzFz7zcg0M7p/UETExIzE+sNC3v9GTExEc9rqdLdtI5LpESCI9n1P1pl8WrCoXC7E6kmROI55PUcmzpmWYR4Uos30U6/w4eM0ep44kNdrr350KaWUUsoPnwqgSymllFJ+OP3O73w1RiMnmAhyvx2f/b2Xf/gzP8PtPDVBIESCmFkYe+9769xVELDJ82rHdZ7PW2+UPq7P5/XJ7eyi60CemfPqKc9pZpEhwsQUPkBgJkpkhLuLKLMk4GbuLqqr5JuRSSAiYiZmYiHwSjZJiIXCLBPcFMwAUUSCQIxweGRGZrr77XYjQERaayvdHnOu2nVmeriNyUTKPMbICCHu+8bMbpaRAETE3MxmU2WicAdARCzMLEQY50hAhIEVfceaUl6J7T01JgJgbp5B6wkwPCIyMrB60DYt1uBIZEYic10gbL3dboe7ETFAEWFz0kq0iSLD3VtrIppIZBKRqgIUgTknM23bzkxIuHtkZAJJrbV9267Xq7mrqqqu1xaYiYXdHQlmAgAiZTYzj2Dm9TnKSIBEJNIjPD3WZnREArRuDkbEnDbMk2jfL5Y5zMHcLpfHN94AN8gO2U+L2zCLuI15O+c55pguDCEFBIe9enG+fPn4oxfb4Z/5sZ9+fHzrL/z8X12PtJRSSiml/KCr7+pKKaWUUn5IvPPOO62FUmwSDcSNrN386VEimMFI4twa9qbgUCEWAaeP05+f3Cd85YwTEW9cLpQxz0OEGaD047iN45YeqtKajjGYuW+buUUEMbfeRGScBwDh1zVlDxImZiKKiARUGzMTMjyAZGaogjnNCEysEF4l65xn2gizjABSiBPIRGZkhJtb+DQ7x6miW+9NlJiS6N6tjshIIiiv4JXtPDNTiHnfmDnnRCYAMMI9zIQFuOfLBPAKpqdlJhER0xwjIpQFKxtNWif/iDiBiBw2E9i2DlrHEs0jE2AWz5xjMouIttZUlIhWXoxc7WJmETOLcGZu2kTV3ZG5uscJWqMcLHx/l0jWx8i8hjvI3SMcmaJNRYVlznm/asgMwHxqU+09gTDzMZhXhs7uHu4kLCJr+gMgFkG4u40xADCzirIwEYEozOM4Euv5sLtNmx6x+tL3CQ7ZLNOSSDfWTro9HyOSWLS15p4fPZ1npjkcRAE97V//j/+T3/i1f/Dq/ZcAqbQv/jtViy6llFJK+QFWAXQppZRSyg+2zPzOd75l5/MH73/36dDHR+8+FE1VWpPWlJhUOOeMcTQJRUac6TNzNmUK8/Nqc4YbgDCHx2W/rC5wZhCRiphNMwszFtEma7FBWg83ZBKz9M7CNsY6IQhiEBK0lqBJZI1ysLy+9RcBgJghAqIwW63iJCRASPhIGz5Opvv4w6oOi0gibc61pOzhIqKi94lpAqsA8AhKCLGqhsecnmuCgwARYubEKmq7W2YykbIgc9oEkpiaNjP7eKpCVMMtPMKj9abakng9FmYBXofRIrrvQGaYm0dmJkg4Em5BzCLSpIkIEZm5R2QGMxMRXj8uEWUmAnk4EVQ0MjIzidaPjAwiZpKPa8Lrf3f3iAAgvFJ8RNynt4mYCBGeRKD7qwDpvlrdbgYQEa0/H6xHmaBEEpDhYwyPAKCqBNznOzLZHMgV+Gd4hHm4r8cUnkTELYmSOEi0b227DEOSSN+lbcQyQjx1gI7bOcYRkWBxIMK39mDjRIzPvH99uJ0/8YdP9OUvfwK/x0oppZRSyp9ABdCllFJKKT9gMvM73/rdcTw9f/geMx7f/JHP/cv/6m/+5te3OM0zPbauD/t+2XoXIkrOQM4Y1/n0IWxSOuBzHOd5PF56V2XKCEeChdMizIEVUfK0CZD2tm7lIQL3S34AEZjhjgwQrSIz1nhxJoghDBGYIQKqiID7GoZ2D7yORe9d2oiIcHd3zwxGIiPDwmbr6zjeut6X+76DyOZY4x3ERESZcR7DwwGwcALuLizKTMnHcd5uN2FaMbG7MVHfdmHOjOM4iLn3bWstM47zBkBYtm2LCDNbGffWNxEJt+vz9eHxcX94AMsYxziOJo1YkrJp495z3ygS4YjIjIxMogTh/s33SnlXrntfWg6/3yZUbapKzOFuc2YGCzdVMwskr/AXmRkEJhJiWmMjK7te6TOACF9DHxGZgcQ6osgEGmOOMVhYVXpTjxhjPD8/t6at9cgwMzdjkQDMbPXZbc45zd1FOMJ9zibSRbvK+rRFOgNMGffXBSwRIIBEVIl5WnDrfd9ZO0uH6DmmBbRftD1w69ebO4hUk+U2/JiTHO6W4I7jr339D3/9L33uwxc7gMz4t/6j//R7/juvlFJKKaX8/1EBdCmllFLKD4ZvvfOOt5mU25svPvsv/Su/+fWvMbswkfDe5OHhYXvobpbzkODMkW5bkwyb52l2kHtn4gzKyPAkSmFx47B0I1WIUGbaDHcmgio1DQ8keAXNHvfNCgDEYIYwfN0bDODelV2Bsk0DoE3X0b1MZCYhicQj3dwzAGLlWKXfVaPNNJtYfd714xOqwszuERnIXLvMmTnGcHcVXVvPayNCRIU5wo/z3Pe99w2ZNs2mb1tfSaibEdHD5YGZIuJ2O4hobTEDMDuRIBHtGwjp4XOQiG4brVrzeWpXVc3McAs3JlnVZSYkcmZK76oaPsd5nse56smEXNXm8HvwTNBMyvsWM60P/N5xdjezaYOZem/neZurdS5CRHOcq0Fu01boHBGrig7cHw4z995temSCaG1kj3HOaW7OwiIsopkr24+V5t975EwsQqDMWK895MdFakJGRvred2GJtdzhnhH7vu37Nm1G+ppLISZtKqJEdI4RCWbp286qmWRu7uGB3vfW9+n35y7bI7NMi3Oet+v1ehyH5UhONCJ2n9w6WD/zYz99eXzrpz7/hVqLLqWUUkr5flbfq5VSSimlfF97993/STwQyRN9buPhSslNmYXCB0eo0MO+aUMAPA/2kzLdhtlkRrrPOeYYjLz0ndbqQiYJQzTPE26cQa2BOXyGO9KZmURSJSLuOxpzwlxY1ggzwCTCTX0aMpQ40iMCGSTCIvM8M1JU1ihEejATsyTIExHrxB3AnHS/6BfIQEbEuuyXkQxqoswMInf/OAFdzefjONysqa795WlzXecT5swcc/Zta71nxOoC923T1wE0g7beQJSRww2ZQgRiIqyslZil9RVtwxxM1BSR6R5m92+iI4BA5us3ygwPN4uQrUtrNsccY45BRBlhNrbeVSTSfXpYimxEAvDrEH4Vmuk+nJE5bBBh29p5Hmv25B5Pm60fP6etJ7YiYLlfGsTrALq5Z2aCWVWZaYzhvj5/REQJfHzVcMW4a9GbVdbJQfzxdkcyC5MAiIyM2PcHEblvoWSu8et968NmZrJQMq35FyJCptk084jc952YbdpKrt1cRFl0DMsEs2z7A4uax7SYAQeN4NPJIAYycCSSCKm/8O/98j/9+j/4w/feO4O+e+1f+lKtRZdSSimlfN+pALqUUkop5ftLZr7/3jeP6/PTB98myrbJVN6mm2ekXZq++akX+95EAtePzucPn5+eLk2RcdyuylDhdfYPyON29fB1X44TXZuNYWMK87rj5+7CdNm3zHSPYecKeVXvmep0y4SI2Bjpcdn3DKxpYxXp+34eBxKPjw9mNubMdFVRbXNOdwfSPcIdEb1vvfcxLUDEcg+jI0gAJs/wcI+QputooZ1GoMvlsmJQD0eCiERFRUXEzTJCWUWEmFamDaBpY5FkWdcIkXlPd4VXpJoWcKe4V4Np64jIcxzHANC3HhEEiOocc8yhoiBEJu6xcK6pkLWrsVLblcrbOCNcREg4gPM8iaBNwuM8bk9Pry7bvvVGTMf1dlzP1i6qm2obY7hZZrIIAXMMYWmtWUxiqIq7A1BV98jMvXdVFZGVPsv9emGIiKqq6jqluD4+4vtqCtE6Fsgr6HZ3MwMgzL13FllB9uuLgp7r/iELEmYuLCoCYH3423ZRUURABMJgRgbcIxNM3ARNQURzut9r9e5u5tu2efjtenWzVZk3izHGq1dPcxqBL5cLiQ73dBBJ2zdqO/rl4c3PBLcPjnGOMDMwbRDAovu7Lx9/YvuwYX76/XO/2U/90XOtRZdSSimlfJ+oALqUUkop5ZOXmR/9s392nOfzB9/dPvXmT3z+537nG//zOaYQ9o0fLn2/NADjdiM/G1NrqWR+ezWO63kcvTUgx3kwrV6yzDGO4xYRzKTaVqLaRMIjI3rryAx34B5QijAR7N4yjoxAJmjNF5O25tPCQ0VIFMzzPJl4u1zcZnowUUbEPa9kBl7Hl5wrB/WQ1ljUxgkQSaN1uM+dhCCUyIjICGqNmEEId4oUJiIGKGlFybkqwJy5pidY9D7tvGq4K3RlIhab08OFVxq/zuRlZq7Lg3OMyABR3/eM9GHmQUTa1D0iPDLXvISqeuRcATFLa30FqeaWSGZu2oA0N0qsSDqQnvG6zU0JZEaECQszZQKZlKzaiTgi17bJemIEZETT1lo75xkZRCTMLPJx0NxaUxEivl9QZBFhgCJD/vcjHu6tNRFJYM7hbiLSmoqqzekRmakiwoLX8fSql4PZxolMESFVgGJOAvF9jiPCQ0Q4AXN8PHCdcR8lcbdwUknA51yvaojINJtjtNYj4na7MZGIbNt2jnkcp/l9fLxpT9A5rLXeWmPVAIfo/uItSLcg6RfRLox0H+fx/PR0tTmnp/AY+Df/4R/9+l98q3k8nPaTf3CrJLqUUkop5ZNVAXQppZRSyicmMz/8o98/z8Nt/vjPfOGbv/qr195bS+FINoAbY+u8d2mSknM8fTiP5/SzCynTGFc3iwwRISDcCWAmbXrcbtfnZ1592NZyVXpFM5OAbdsoEeH3cjGgykQU4QCQ4WbIZAYAYhbVvO8sJLfGrc/bjYC278gMMx8Da79YldYixlqLZl7d23QnEbBgDoBIJEkAUASYku+7E8hIFjAREzIzLMYkFmIOogyHO8DICLd10C9FEEHu9wzb12gIich5O+YYoqzMTGRzunlmCjMixxyRScytNSQikkhWBhuZFjHnBJKIhMUjzumrFr31PUAWMc8zARLZ+gaCuzHLuojoGYkkZiQyAwRWab3hfmsxm2rXLqoRaXOu3YyFiHhtiYiec6xP8bb2Q4juTWdVYSbQnDMymKhvG7PMjz8RzOuCYuudmTNjjNNsMlNTERWbtl5d6K0xsdv6V4gqCYPIxkh3Zk4RALS2PNYKCogBRKQ55szw+wh4RoRb+JjzHCerEtEfj0cLe4S7t7Zl5Hkeqtp7v1wezjGOc4iKiLIKgSJyTN+2vfUtkJ4ZgPYLixKo9721LtIyMc1vt+OY/jzPp9uwwEwhCW7+13/tu7/xs2+90g4TvdIXf+VXvme/tUsppZRSyscqgC6llFJK+V77xje+wXFK+ovHh5/42S/8/j/6H436aug24heP7WGTRhHu4/Z8XF/Z+SQUD7vO47DzyJh719Z0nFci2rYtIojRtCETSGaKzFjn45hJGOYAqPV0T3eRBhDCIxxMpJJxP3rHzMIcbgysJYfMzAiWdp/yYGbV+5A0M4jCw8dg5jUfAdwHjTMiX7eOI4KYmHhFvAA8IkEifM8n72+YZg5KESYidztuxz2KHeeKYok43OccRExEkStwhrKExxhGTKLaez9vt/M80631trU+zrFK3701Xb1pZhCmGTO31ps0ADZNewPROYYwa1MCEhQgXYPUYNp2iMRxgJhU0xwEFgGQGZkOUVIFUbqnm7uRaLvsMEtbKxpJwFq9yMhpcw2brOXlfD3AvFrYNufDw0Wb2rQkrOKwMBMw54zIFUAT0XE7ATCzNmXiBERlvxEAACAASURBVO4b3BGvF57d3TJcW1vF51UQdzMPjwgCsTAzR+ac8zxPM0ugN3UPcwOgLE0158wxfVrGyofhbuaTmDxiztm3rW9b7909pllEtta2y771nYjmXHXs1rfu5vesXAUsCM/ITOLWkthWh5oJECSARBKSABpjHMc5pknf+uXhOv0IvBru4KSURIR59u0l55vXlAlKzvzil/7z793v9lJKKaWUP/cqgC6llFJK+R7Jr3zlwx99cfbt6a23brQ3+6gBLHh86NrV55w+yb1zdspGnu7juB63J4rZGu8Pm48RNhGmIiJs58HCul/SBjJUJd3h90mEBNwzABCFWyZIW7pnpEiLWGFisrA0zcwIN7OVfK4ytdxXH0SYV5CMdTkQ5DYjEq/jyxXsMnPvPSPMLNc+BjGrENGqVAPIuIer0y0BVSVgrSoDyMzjODJDVVtrEfH8/Ny3rfdtjLFmPV5no4OZiXmVcYlIWSJyTidmEdGmbuZmhGyttdbGcSZStcmKrkHUlETMjCIYqapE7JkMEOCZpCqicAcRRCmCVpm3NQin3TdMfFoiwWxmGU4EECXgsU4Urgg+PddZPkJSRKxQXkREJeIe1xOzCEtrRJSgDF8vDQgTEGa2Ku0EXjXxtbWdmcKCxBiWmbjn1wR6vYVCJEygdLf7vkrS/c8CFMgIj4xcxwk/3or2iDHnOEcCj4+P0+0cIzNFtLcGj4xYByXXWUIWFhEPy/WpF1bVvvV1oZGIRURVhJWYk8AAA0CCGCC4rV83Y0X06QFzH+cAEkRuq7POcxqA3jePNHcz19bavp0J5x7tQXRjVs5xXJ/GOOb00yTYNGICORo5t+OhOtGllFJKKd8D+km/A6WUUkopP+TeeeedhikZ3zyPn/zWd37/595A4i0dQaoConjYITiNXqkfbiMsfNWE09OG4ty6tq1pVwhgjGzrZ+ZoYCERckZ6+EwzmK/NhySMc3pEEq30eK1hAFBp5n6OIeuunOu9leyWkbkGNBIAtt63Tirq85xziggSET7WjcGEiqz5iHAHgYnS/Txu7sHMvTeSDcS55jUi10aEiAyzzHRdA8R5nicAgK7PT2vj+HK5ALA5Rdv9WiALASqSSNAKOEW0AwCSIAC1BF7PGbeNhNfRQmHm8xzEtO37qoFnJPUO1R6Rc8Y4RZiEmSnnhEdThTawYEwwQTXPI8xBTHbCKImApAg38wjPmHNmhgiHu01zs3U1UZjntOvzc9/21joTeUS4g0ibtm1jEiaie7xNTYhEkBSR4aEs87yZzXBX2kjgFkmUxGHDzdxtrFQ5ct1KNJsRuTrUa9CDhdayNhMReIwZniBEzAzLSCJmFhWNzAjX1ohlvTiw4myGEElmrD44RElo9b450+bc9v1yuZznSUxb3zyMCK01Xq1tVVpleA8wta2lWcw5z8HaRNSOAxEivOazV416jjnGBEAEm57EIm2ME0T5+IaoqjAxsyTBFClIZSh7175ps/54u+mHT8/I4YALpcP6+fD+Z277q//mK/9liJ69/82/WUl0KaWUUsqflWpAl1JKKaX8mfhf3/kqiInIoc/RH3DtCWhrXd58fNg7n7dn2EFxIwxlVwkIAYQAWZC520Q4EMggAjGHjXsAuq7teURGItMt0jKCKRlYDWJtepynhwPUHx5F1ceklduK5NqAZgZh1YrXz+pm7q6qCYQHrSovcs7p5vfiMACmjDQ3Yab7IHBkBtH9Qt3q0rLcjxCut2UiNyeCKnvk2lkQESZy93U6cNokUG9t2zYR8XDWxqqZgdXAfj0qDRESJWkreYUHWNDamqWet5u2pq2RMCUQSLrH1qvw69N8Ze2RTBDmtX49xrk6wmv8mljCbEXeNmeYeSQByJxzqmpTdfdpNufsTUWFiFYxWV8vjqgKMyOz901E1yZGAtIaizCTm4MgquZuvjY61nx0eNiqcmc6r4nqiOv1BnDTlmtVw2YGmKW3xiJIHMeREcIcmauZfr9NCFp95UwiYmUZ42Y+M1y4tda3fQ/38+NNlbXizUS8snxlZhAl0iyIaOub7BuYx/MzEzVt67ULAplPImzbluE2h5kTkTKf5xmZouI2bc55nsikBJkzk6qYubuvcXNmIcJ6TWHvGzGHI8ITYBFpKq2RrldQMtc8tch5O3xOZblH8tzQmki/jfHB09OH13kbFCIk/aMXL16MYw2yoMm//R/8Z5/gfzRKKaWUUn4oVQBdSimllPKn6d13/z7sgYIxxW2AVYQ50YVXV7gJP/Qm5LdX3+Y4VSLsQA6mIGEAbsEBzgzztYxwH69YUTFAWIViNNVItzm4CTFlOK/BB4KqqMp08whKtN6ZJdbCBrD+lvejcpmRzATi17vQAWaAIpJAwOqjri41rWS0dQXIze55MJBr/jhirSWsqBREq8q6gmYVCV8/ACDKTA+X9VzWbgU4AV4bGkS8YveMSDDdVyVeL0iAREBsATcLM0IyCzWN8JgW5ylNWXS6I9cYiEbEOIe8Xl72cI9YW8mZqSIRvgLodY5vndUDVt6PzCQQM88xbBoRNVVt7fXMBXrvIhwRkQCREq+nrF1FRYiEeCXXa607iRKIjHRfLe91pm96AOvpuUW4OUDMpE0iwszNnIhZmgiIgAz3QKK31lRZdJXZKTMimKWv3ncGE98z5SQmFhbz4T4znFlVWtu2iLA5geT7PURZKy4iqk2ZORNx/xVTiKR3EN2enpApLMRYcyJzjkCqKhMi/HY73WwNfaypDREBweaEJwEqa/tkvRyyPmO6Xp9YX1Fb6wTEtPXF5m4szMKr4x/hYZEgFrY53Szd14FEAosqazuczqCnEYflgDhJiKYIO+VDb+Zxnu5u5+2X/s6XP7H/iJRSSiml/HCpALqUUkop5U/BN77xVXGiJOagy42OH2VEhmegNWqUG1xzCFkjiArCrh+9r432S89xm8f1PJ4JEe7jOFW1tQ7QnPOcQ7STSIJFG6siyS2QePPNF0Aex21/80XbOhAYE+5QXgkzhICEZ5wH3Jkl3cMs/X4e0N0Rec+QVwIMyqQxLQBmVVViDiS9Ph5oZm627Tszf3xjEMBKnF8Xn2ldEQQQiUgA0KaiDa+v6okIiDxjxc3UGiLhSb2BGRlxHHAj4XmeNmcTEWEQbIyM+1tF4HY9zuOwOUVZmJQx5swIZWZm93j16plF+rZra+eYH3zw4X659G1TaWuhubftHON2u10eHkTE3SOcmfq2nedxnjdVBXC/obftD5eHDz/48LjdXrx4oapE5OG99cfHR2LKyDmn9k1bh/kKkGXvxISImMPGOI+DkMg4zmPOaebCHBHHeYB53TlkVVYxD/P0IGlde+u9uVtkXi6PzBIgbdJUtqbnGGvMuvfe+9b6hswcw93B0i6Xcb3acRCT7pe27TEnJVgFlEjHirzBKQIiQsIMbomEMoCck5CgVcxORBIj5hzXZyJy9+v1CkBE1syGmY31sbnvD7u2frvenp6en6/XFy/e0L6B+I0339wul/AASES2bTP3Y5wvXjxeLpe27R+/TnL/+oyEOcYJonCf522daTzP0908/LyNTKjq5XJh4eN6dbf/jb23+ZFtO8/7nvdjrbWrus/XvaQMSVQAB0GEjAwEHimZOIARQ0AmGXCWTDLwzAMjQTLkP5MJJx4ECBIgCIHECGyAQRCEtuJYhhybImVR995zTndV7bXW+5HBqr6XpCg5SgBSlPYPjb59T39U1a46hTrPfvr3hLvPkQkQjz6mI6XowzvaHkwrnx5DeO8WIPL0yNvHz/XUjCgpHfQ3j8XCg4ODg4ODg4P/fxwB9MHBwcHBwcHB/0fy29/+0evXs/HzY+MaXdCGBIGFTyqvzxszIYxspxgSE25IozR3DzOfOyGY0mcPnwivVZXJzViERcF0X67TBtFkZi0AZ58JELGu7mv4Ws0jQiy78Wq3Uu77DmQtJcbMiLuE1+/2YWZenWgVIQIBYIZoioY5QGDhFSKbUa1UKwixd993LYVVILJm6LC+l1f9Ogl5d3UQh1t6IJNVuSgSPuccnUVYlYrenR6gJfxVLci0OcNmZjDTnNPNquqSMfT9lhEiuoTUc97zdCCZUgiRQQQV7XvvfXhkqbXWbZpZRGa27UTEvfe2ndq2Le/HmPN8PjPzNGMiolXj9USoamaaWd22UquyzGkeqa1RJuYcYzDztm0RMW323leYGxZEYCEWiYw55hy722RhAgjLl5LILEVZGKvnDLIMrVVbXWYRc0ipzKsWb5morTErwLhXqN3NYuXyzEwcHsxcRNxWK/huGJljgohEMoIAZom0RArW5mF65HJ5r9uPDDBFht870S+LihGETLc5+hKZfDkjGRErTV5nOPoYpdbWmoquzUApRUSJZO1RrtlFEdVaiCgyALoX84UJZG42p81JEZTJGZnwsDn2dM/0iLj/agCxsLBwRLh77/s6IGEG5PKJAJTg9vio50fUjbYHbg9OEoE+5tPz5bmP65hE1sHF4E4eSOL/8D/9L35xTzYHBwcHBwcHB7/EHAH0wcHBwcHBwcGfme9973tq/eF6+cb3/+Aff+MbrXVwllKKKogZJLAzu8IoLeeePpHGRMg14DfTXISQke7uEwRRaUVVCJm4p7dYS4ApJYkjAdEEqNv6gpgTCWKaNiOC7+ttnpEsJEx935FZSrlrK4iYmInWMB2LhJsARZWWcDgTWkgV5iBmubsXbN9526RtxBS9++0GIlaVVtMcGUQEplx+jEhkLA1wEsM9zcyNVWVVic1sTmYhFSoFS9yRNOacYxTR9Ji9R0YCzLQUHrXoiiNH75mxNBpMhMzla4gMyqDlNhbmUvbb3sdgkaJFWfu0ZNZaikhG3va+nU7btmWEu3t4a42Y3YxZANicRCBhYc5M81h9cMrE3YNMYeZ9zNETUNHIVbedHrEOOYuICgD36GN4GJClrH42NxECMqNWXZ7o+xpkOhfVUgByzzFDRImWUSMyE7TU2xxukb4sKflldpyYY6wU2N3d3NyLKBPGGBkBIO5akXvx/UWskcvUzMzhHr683gTAw+KeO98zaF6Tgu4rei6lLEOLu6nq6XS+GzY8iFhVz6eTqCZo+adJdPTd3VWUlpNjHQGm0cdYhe51W2zOOcxmTCNg3R2ZGWlfXkNmFtFta6qFmcaYw6aHl1JLKemGDM6sL76XUouWmizQitKCJKmA23XE8+32/vJkc1rQdOwTQdI4+BykZK/2v/E3vvULeuI5ODg4ODg4OPil5AigDw4ODg4ODg7+35Lf/vbnn557kafXr6e+2fpH4nBPZi+cb161pqyI9On9tn/8Im1QrrE9y4zT6cRCNkdEMtFp25iZgIxEUTqfyAbCwYRwuCMCd1dGTPM5ZmauLA+R7h7uCSIWD08i0eIZEQEiFhbVwrKqu1IUwOhDi5ZWmXk1nsONKatqeoTN0XciIuK1X1dKAZPNcXt+0lJKqSycsabjBrOctlOEIyEqmeHh4b6ECXfzM1JYwv16vUqRWsuyKQDERAFYhLllpIhERngUlnSfc8aLKJiYmEXXXh9JfKVkSGZU5TXll0npkdN5CT3algggwYxpOQy1kSpEaHZEpCghKSPXoQ4nlmWmXtl/hoMELBQBoiSet9vdo83ITJtzjjHHzLsnO5iZWZg4iJKZWUmEWCzCItyjnTZVjcwiWkqpwuk2xq4q6/wEEKDkVTr2EOE57XK9ESCqp21jonDfb93cM+A2Rai1hlz3oYNAROnJwlrUI+acvY+V1687noB4GU7c2klV8SIat3UrhPd9TJvhKVpWOD7GGH0Qy4qkWdfjl8wmEb15/Wa5SjycAGaurdXWSjvZmGGz1soiAOAOAoSj7+nGLNb7HB13dzhut91sZuYaKbSlGme63W6ZUC0JsHCtNXG3vqiW2ur5fC6lELNHJhGLaKtSCzJzzhhdMokZVWn0HMM8wJIsnokkgPswJ9bt1C0ut/6jD5celGAobzjffvW9fjzfxitDec7X3/zmN38Rz0MHBwcHBwcHB79kHAH0wcHBwcHBwcG/nu997zuS8XCx3/gXH373N7+eM6WUU5FaCnzCJmMqh3AIQhgUPvcr3IFIJCiTUFgI6TaXL4NBK7UMDwhzLT67zWFuRbWIZni6RzgBmYhIomRiEaEEMkAMUCYgDCYi9ohA4GXhTbVGxNj3UiuAW9+JaQkP7pYDd85kAiLCffSdiYQZGUJrIy7dbfZOzEy01vYikwjCUkTnHBEhKkSETHdbrdrwiPDILKUQ0PddhEspxBQRbiEixBRMa7FPi4a7m1cWYSWRFTIzEYhJmKUAQESAQMyqFIZwprgbS8Dp6dOJKYmTGQIiZCLMYnrQMj2Ijx62JCPJwHoDcrrf+8WLTJAQMb0koz6nzenuZhOIVhsSET7n/dwAkAAxMYmQqNbKoiC2iMgMoNTKoqsdTURbKUwIN7MZ6UKUGbgXx83ciMg9Zp+ZCYIwrQFGAG5hw0HBRLo0zYnVjWbm8NCi7bTt+z7G8MiiqkuZkoHEywglhAVJ5q4qLOz3AcU1zHg/DMxSa70f/lzSFAIBTCzi7kR0fnwkQrrfe9DmWlS1iOgcw+Zcvpj7TCUyM2bfYw56ma909wyPCCJej3N3c3cQlVJLq060HhLmQYTa6pJRS22iKqIqtEwjkUggmcG8dg5n3+ftGvPudeEMmO17X03z275noLC6exBxLQZ10uRTlOaJQM6EJRwSRH/gv/51/EHx57mPY67w4ODg4ODg4OBP5wigDw4ODg4ODg7+RL73ve9JXAhO6JNRw4mkUGFGSalKjZ3mlXISlq45GanCQplhyCAABGICs8+R5oQAcSZ8mpt5RJiDIMo2x5xzzNFa21pLRLiHO4sw86qv8ssaIIOWKSIzSRSMREZG3vUXS3LQImLsN9UCYB89V7+XGUAAFIkMhGMNx80py5nrxkTCkhmr2rwuaLWwQVRKUWEG7ftu7qososQUHuvC7yuH4bU1YfE5iMAsLOQeNqYWFVVSDoCISinubmMWllJqbacVHoc7EUOEWO7bdh4Q0dZgM22mTyIilkwOD/8yAA1fx2vpkVe2zExFda4c2SYzi7CyiAgTbqOb+YuXArjnzkwgolUshnuM0XvvQL55/bqoZmbvPRNadAmdAbCISCmtrSTXI5IAXt4MWrcjI7baRJiA2351N3454EBamIVhqUwCACLCfGYEE29tc8/Zp+pLiz6TmEjuHo+MKK2ezufr5TLnZJFaqojcLeERBIiwqIaTe0ybtRSt6svonCh3UzPbnEi01lQKMZsZEszsESuAjgiApLUMjzmZ2d1G7yxCoIxwczNzm7EuerlE3Kx3t7kEIMQUL3fVtp1ba6XUSAdSRGvb2naSrRILMucYmSkiZkvGfSIRgCgsbFjfPWKVySMRmaP3MXbr++w95oC7KlPmvndtpbb2/PwMz6aFmBJsGcnMWtv5jbYH2c5yPnenj/sckVjGGczLF0/14UTCSfj3/uPDEH1wcHBwcHBw8LM5AuiDg4ODg4ODg5/B7/zD/4FESevU181/lMSEKJynTRuDlhY5Q1b5mJmVWYQBZKRNtzHHjnQmMEiIiPD09ORm29Zi2ZYTzCwiEUFEqpoZoCQRICnBKmvTjeTeL6YMZGQGgQmUdvcteBjSV6oc4R7mvkzQClDm6pXmMifkKpwCAC/VRIatQnR4qhZhenp+BtC27a5HjiBhWuKJ9QqSSERKKft+c3dVFRFmYRFaUfldY4FaC/MSd0xzY1pJeaiqqNybzkyiisx0Tw8ChIVEI3Jer0QkIqyKTDe73q4eoaUICJEZMyLX6NwKOrUUJnK3tW5oti555fjCwtMs3OkeE4uqqqqwjjEiAsxfdqDXDTEzIJmptsZEc84Vc9dal4p6SZCZWIsycYQDSaCqxd3HHFizkCw2p5m5OQG0WvCEJLi7RUSkL+VKZiBXB5lFam0qJYE5+1Jat7aFp03fTlWYI8xtJlJU162mTFWtta7rpqJfJuM+bfYOhIiUWokLQBmxuuZZBBkwp1IgAmaMmWZkTiwArs8fKbPVZr4k3WxmZu4RhKTMPsbovY9dVTMxel9HA0QirKIJRLhNE76X0pMpCaUWYkai1lpr27YtViGaWVVFC/HayWTfu49hc9wu177vL0qZVMKc+/XyNG16JLFqqVKqWzCTKoeZjd73610bzSJVWXXOmR6cfDqfAvjw9Kytte1E2kgqSZlBqJu0s7RGWj3m9bpf9uk2g0Hdfc+MZMi//5/9lz/nJ6uDg4ODg4ODgz/nHAH0wcHBwcHBwcFXfPe73200lb3QnN2lnkpFFdbCDOfoiq5p4hbuGUnJUiqLEBOXkhG+33wOt5kwZBKSE4ykzGFzFUvzRX+wis0v0gNixlJkLEMCgPAIdxJOZLivSrUIxyo6exIShEwPN/dOlLx6w+ERwayEFUtnZvIy7BIi4sueLhFAd99yJrRUVrk9P4OotOZmkUkid3syXmwgESs9tzkjk1UZxESkSkRrCXDN2/G9jU2j9zm6sKy9Q2EGcwKea15RKZHuNkdGMhGxuMe4XZmYmVdMT4R93yNCVnhMTAh3N/Nwy0wmqq0RcE+TiVTVzMaYyw68MlNmQhKtKUBetW+OXPIJecmf76+V52rpqqgwgSIil2aDeWlDVNdC4OrGIjMRvpwScVd1B5BIpHu425zr+gNrcJKTKJZ/WYRYIpOEWSSS1t5gayciGmPXWkqtIiU93b22yoTwGRlArgN1v3dYhHmdiqD7rWYiiohwRzoyQVBtAM85CUlCUIlwH9Myl45EMsnd+linH9JG+vrM3fTi7nNa752JVXj0HhHEYGYA7i7MRGRua36wtY0IY4xWW61Naw2iBNYIITPT2m5U/fLMQuQqZgcRkbLt+9z7nHPuu83BL78ToMpu43p7jvBMMKvWpqUSiYjck3qfc3RmVtW2bXxfSnRKUpJ2OgXw8fm51FZbAyuREIlFQouezsRCWiDFPK63y/PzbZ++X30OkyzJY5hm6tjbb/+dv/MLeAo7ODg4ODg4OPjzxxFAHxwcHBwcHBwgM3/0g/97jucP7z+/+vkNX6WacCEmkbIVnNkxn8guFFOQDCISn5FBXDdiTiSV4nPuH967TyC0KDKRQZmIQEbdmoiu4A6J8AASFO7uHp6x2sOZEBEmmjZtTDNj5gg3myAIS23VLGyakBDlctq6jev1SZhURZhWxs0sACNXJxZIkDAzL40zklRVlJfomMEgSK1cSvQOgEXdLImkNSoFKojMCLjDV3zJyAQome8GYmHKhPtSR4Ap58xIVp2jW+8qgqSMAFFkWvqYMyLWfl169Hu+zASEx5hzLd3t+y4irVa3u8ahlKKqwuxmZpbhKlJrba1l5u12W4fu1evXbtZ7XyJsizidtqLlHjeDMmklzqKFWUAEIhAy814QjyAmKpJmiACYVEkEQL9e++12enhYReA5Z3gIc7qbzev1SkgViQh3C5tMRIn0WH7kzCBi1sLCCTKPdjqV2iJDS9FWI2GWc/p2OjFz36/aqtaGBCIQmcyZET6ZiQjLbOEeKspEyJz3zrVtrRUtYUbCrIwIs9F7r2VD0u12IwILkdA06/sco8853awVZSIb020i47yd3Oxyva7muJaySv+3fVeRUmqYlaLnh9M6HyCqRQWE6/XSe3f3t2/ficrofdvO2+nErS4tiUesYnLYStEjER7eF2NkJhGUed/3OYa7UwYBTMTEQqxFEjHnzgyi9YsJKlpqbUQUvjw5AQpVLaWcthOYItMthLlqlaIBjDFXOX45b5goiSGKUpYHfC5ZOItofb7290+Xj9fpHuagUp6/eHV+tUuFFP2tb/7dX9jz2sHBwcHBwcHBnw+OAPrg4ODg4ODgLzX/59//+6T28Pbtr//mX/ud//V/1joLsxK0YCtVmci6wiXNx5UyVGgFyjkGkjIxhyUCAi3F3W7Pz0JgJiIyM3erS6ABiAoxLyltBGJZFihFZO2wuc9ECjMxEygzzNxsLhnDfX9NSFjd0zyZVEsptbjNSAfgbhmhKmv8LWI1bBlERFjLbiSSa8CQmQgkhKJkAzYpAusLzBC+urLhbuFFCrP4tFVIxb3QC2bJxHTzcCC1VSJCfOWQgHtGAFh9cCTdXQwkIA7K2+02zGqtq717vV6I6LSdVltWRCLjLimu7Xw6r/SPiIoWUWHmteW4DCGIWKuB69uJWYtmIjKYKDLd3cwIqLWtvTqbZu6RUesG0Jhj6afNnJmK6HbazPx6u95X+YgSIOaiOuYYvRetCdi0u5qjbXPamNPDtZRWW7gjkwlzDGF59+6diGTGvncmKq1FrEQziRlEQK5TBW6RmQRWFne/Xi+Bey5eS6m1Xi7X3nczq1WBvF2vRMwk4b7iWmbJTLN52rZWNMZkgggTk5n1MVZBfYmbM0NKNY8xbNvO5vbxw/tTa1trW62323W/3drWhO9ia9D98BJoPeRERFlURFWZmQgZLirM5OYRlpnl8YzMebmUWrU1qs1Ht9vN5jCzMFcpGdl7NzcPn2bLKVNbYxEiMlunbJbt/N5hX31sZoCibZuqujuzCAurZKR7EIKJVjmcCBkpzCyyNiGZ2MwSKVqQmeY+OiNF2GxpbBB+r3/f9n3vPSFaz1q26ehuV8s9wiGBWk4tM7qyE81Nfvu3j0L0wcHBwcHBwV9SjgD64ODg4ODg4C8jmd/6/Pv/1pzn58//iu0pW69bbcpaVQQUM/1Zc5Z0uS8G+uwdmSISbmkOs2Vj6LcbGFqVGOHW9/7lVOCa4WNey3Cy3MkJJCgJWDZlgjATEhlzJYAs60oSv+ib3YiwhBN3F3RSLuWAqtZic2ZCVTwyMpnvaaD7Um2s2UIsjwSYMyKJkijTk5DCmB2z++gswiLWO0UIwdw8jCKVhBOzj/UDk+4WEZUCQp/Tw0Fop7ZuOCGRsORMzQAAIABJREFUmW5rdy/MV7HYLZYYAWuODznn9IxSGwgeMc2IqJWWSGapra3I2DNKqbU18wCwUnuAwMTEtHJHszlmIgHIS5c5M+ec02atdX08xojIJd1e4fgSPRBJZtqcy6cxzVSk1XY+n+ecT09Pd3UJU0aAaWtbIt09AxHh5hHBwnU7TYtp5pnLZWxzElC03G5XAO/evSPiZeeIyESqMACPGL17eK2FCJHp0xApRGG+LNfmnpmidD5tp9Pp/Rfv933PTGHKzN531VJLjUh3c/fHx0dVnXO2qkI0btfCXEuZNiPBwh6egKqYW4SzFBADsp3Obv7x6cOpbadtO21t3/d9v7XWRIWIl8eaiTJBxK1WIiGi2poQI4JZgAybkUFIUV3jgy7k7r7fYnlhavPefb+5WZiHRy01I/d9z7uiBEkEptIaEUXmsp0wCfEStCjx+liYiYXq1kRk9B33hJozERGIICxLdkbGHFOYVORewXYPN4C0lHSPOaPvlMFEY8yINbCJTHj4GHPO4ebK2uoWJKGb15NpneCR6VQcac6XN+X1fi0xpflf/4++9XN+rjs4ODg4ODg4+IWjv+grcHBwcHBwcHDwc+Uf/S//nYh8/598/MZv/h+/+w//ljyMbavM8lDLqeSpGGJPumZcxn716aWeOZDTs3d3N6DvPSNKKYg0s77vtZXadI7pbpRh5hGxNvpKqWMOTpRSlgNXmEWFRZmZhJMobS79AKusUcEVdIqwsDCzzQGklrJWAMOdqLAUkABApoDXpCFOFapwX3JhlsjIFZzlsug6sJwfvqwQ7umRQWFhY79eqmoRff74QZgfzg+X/ZqUD6eTxYzpY99VSmtbLDy4Ln3HvYtaWFaqW4sic5ptrRYRGxPhkZ5IZhTVSHiEm7VaS61SyjSfZq/evCXiOQxgUdVt82Fsk4QTcICKiGottY8+54zgWlupzc1mzEGM1YwNXrfdI95/eP749PHdu0+Y+Xq9ElNG9HEJD2Y6PzwwiTtut5uby5qTTMzppepGcru4WexTRjd3B1FkMPMpopbKsvW5u2W6ZBIlz8FBYqxj2jCZk/cdBJwaXyePMT67/lF4EPD48Nh7f//+/du3r0vRPsbHD+/n6O/evSGiOafNAXfK2C9XSjw+PiCTCA/nTZgJ1Ptuc6pq33uYi0hhraW2Wuccl+vl7ZvXp9PJzAjpc/h+a609Pjx89tlnIvLuk0/Mprs5cs0fRmbbzufTo3m6++m8tVJLKcx0ejhnZq0Vy+x8OrFwukXcHdcRAaSeTpTI3pfqHMDofc7x8PhASBvjcr2aGyifn59776WUjMwIXv18ZvOeme5eam2tlValKIsEcC+wM6loaxuLsjCIWFRU7+daiCDwcHdx88wAmJmYxSfcptlcZhJzo/sWJ+act9utlHK3gbtTOLsjPNznHERUSl2umOv1WlRbKZGM8Nif+zRLDq28nbdX7z795Fe6yNNt7/tsl2vMkFc+L+V3/qe/9/D6V37jr/3WOid0cHBwcHBwcPCXgeN1z8HBwcHBwcFfCr7zne+82rIoHgr6dbRWSaQqP5y2qszpQsF24/G8Xz+E7yoRc4Y5pyIIkR7ukZaxUjIi1lKEZbozcyka4UREpWRmRhBiDdwFgkDClG7rz+9bgIQMT5/AGhSEJ1a7c033uZuqttZoTRQK46VWjGRKcg8i5qLpnuZhZuGRKZQgJJDIZTAQEQBmHi+V6OURISYQgBRhZMy+11Kq1v12ZZa2bZZBTLVWiszpo3ctpW5bZoRZzKm1ElPYfdFOhN19ztlKAXL0LixMSPNlFpkWEObSWDVB05zX4FzbzH2MCWZmFS4e8Ezz1bROC7/ebpfrpW5nUc3ML96///B8HQZiYdHM3Pf9+fl5LqeGx5w255hzfvjw9PR0eXz1SkTMfZmdzXwZM87nMxHZnM+X5/CopRAREh5OROscQALu4WbT5phTVEop27atAzvGWIFyRhKTqJLwGjwEgIS5M6gW7X2YmTBvW9u2TYTXVuGnn3xyOm/IbK0+nE9v3r7eb/vl+alVfTi1Vw9bzFlE3rx+HW4IP29bUabM2+VKyPN2WmcTIqMULUUjIsLipUw9baoKg/reW22n7TTnAEiLAgBlrn8WECVBpKiW9YgP9yVBFpb7cqbICqs9g4hUeJ16UZY5Rx8dACEZmHOGpzCvBvqX//TwWNuKYm7L4yEsIkWkaCmi6yoBQC2laLlby9ejNMJsMpGolNYoA27rDM26E9c5HmKMOT68/xCR93FPYmA97N3NItdftS9TdxCLqIooiCJSRYRo9D3M168yaCnnh3MCEWHTaSk/iItoU731HglpG5cqtUk78+lMpVr69fny9PzhcvWru3j7rf/kP/8f/5v/+vf+5b/8/o/6t771rZ/js+DBwcHBwcHBwS+GI4A+ODg4ODg4+AvO733nO1nzBvzhoF97Fyq8lUZFC0goSk7NodEzLMYtr8+Xjx/ce23KAAJpoCQws2oAM6JsmxQNUG1NSw0AABEhkpi5tpVrIXx9AkQZEW7kTuFIAxIIINJnuoGQxAEOogRlEjMT0Zgmwq3WJeWI9MxEJmcgEp6zD2KSWhGeZmk2RzebzOtyAYaljzlqratWvKI2UQVRBqQoCRNBRQlwG8paRM2dWLTUlKU4YHiE2RyDVUurANJmjM61EPFaGkwkEYW5mReVzJw274t+kWuyzjMC5MKqBSzm6R6RCJK+j9u+J4hYhevltl9v/XrbM5GZfY6PT08fnj6eHx5AMvr40Rfvv/h4uU34i2ak7/vT5TLmnGZuPufybczrdb/d9lo3Fln+BeQq3QaA1hoAM7tdrxlZS0lgZf2rwnuXSoOQMW3uvZdSaq16j6pzmiGTgVzGCCFZmmGhiLBpAIhYmd0sIoTl4eF0Pp/8LrPWN29en7YTM799+/rt29fn8/l2vT4/PT0+bO/enL/+6SvOqEUez+f04MxXD+emKgzro4q8enwgEJBEqUVUxHwIU6lqdz94alFh8ZkiUksVFUS6zbsfXGiJxpk5IiOck8LDbBm3uWp195dCMTHQR0dmq2WMbnMoi7uN2efohFSVOS0ii0iCI3P0ca8ql8KqIGYVIg6QaFFtIipaWCWRtM5LiDAo3Mfoc4yiQgi3yUgSlqLkFmPvt2uGM3K/3TKiFomMOefT8wUgZjGPJVAXvQvZQUQAMZuZmUVkrdvD4ytWAXFE1lpFZO/d7f73rtR6fnx0ZOQynCcSwlJEi6iZJSAvjexEkggrB9MM9H1+9vH2vI89yCP7dv4H//jjv/tXzp+21ub21//23/55Py0eHBwcHBwcHPwcOQLog4ODg4ODg7+w/O7//t9nCBvxM+djukREvHl9fji3psRwH7fbF5/BB4XNcYvR89b77RoRpUmtRVnJISylVnk4s5aMJGWIQoVARJT8kmmapcdaDvQ1u0eERGTaHLPvkpAMSksEMhLBQixkkSAmLaVWrVWkYLlvRSI85sgIm7P3PTMAFFHOhMfoPSMIQKYIt1JWmuYx7+LpKoEYc5xPZ5Uy52RmkSK1ECgjqVYs70ckPGAzPZAAC7GAxQgOIMnH9DnCHJTLZoBwn0NUE5i9mzuAUgqBEMhEIiNTpYpoJkopqiVBM2OEJ1GAk6T3cXm+ffb5+8++eP/x6Xk7P0Tgctl/8MM//KPPvni+Xkcfc9qwcet973vdNrd4er5eu197XiYil0wbkWlryw9Lsp0ZGYnMXDXzACXA9y8G7uYQWh+tgylEDiSgCSJae5IeOSOWacQzVyc9V4j58icKrLMRTJQACCsUxv2y7vK7F38xMfMSgTPAwiBOoAjrak9HZERVfvNKP/1aE0oGEFFZH9r29U/fff1rn3767h2FNy2PDw+t1tNWH86n1mqtqkqnh+3V44OFFZVXrx6Xrtq6L1FGkYKMsGk2E1FEpg2zWbSMvu/Xa601I2/7DQnV8vDw2Pf9ernMMVmk1jb6yIyiEj7dLMNqq63V235DhAqv8yiZ1NqmWswMxKqlnU6iGoCosiqJEgnAABJ0P4ZMstTM7vvtdn2+XK8XQiA9wta5AWRSevi4XS+UKcy36wXprZZpM5O27cSsAN32PTKZ9XQ6bdu2bds6LaIqZtb7cPda2+Pjay1VVImYhcGcRJlYsh1iLm1DUYgCSHdMD/fR++j9fDoT0X69ZiZxCvPeb9frxcw8wpPb+R3X8yD6/LYPSwsilleXt9fH2xA3pr/1zb/783liPDg4ODg4ODj4OXME0AcHBwcHBwd/0chvf/uLr52s1uurahhpVRmnE1cVZLAP8j2jU6bbvD0/MXL5MSRRmSMihbkVZTBAQWuXjwl3cUZEZlh4rtix1Igwm7msyu4JAjGJuMc0N3cgmYgjhCBMAIiJhVWF5T4JuFwPAMzNprkHiJjAyMx0m2P2TDCRqmZEejAxAATAJMwqukqsxEwEpmTlpDS32ioTW+8MYqYVehKQzBHpNoUZEWPvyx2dIAcZyIk8EZFCoEw3Y6aiIqIR3kdXLSJM4C+n4bRULZuNOadPj0wCiZY2pl0utx999tnzbe9uT5frPmaCb7f9/fvLD3742cePz7c+Sm2R2fv8+PR8ud7GmObu7hY+3c1dVD2i92kBc4xA5o/d++s/9NXL3LX1eLeO5Pok8BPf9BUrUE5g5dRrTHKl1ffc+f7Zu+RkRdfrR/Gf8pj8k7+AXt6t2jX95At0YWwbP76SFeeHhRCXUl6dTo8P58fzmTOLcC21irSiWyu1Sa2syg+PpzdvXmvh1ur5fGpVT629e/0W4Tb7adu2WlsRSlemrRa3YXOErZ6+h391ZPPHkvo55+rR19JEFHRvkyOztlJbNZsEqkWJ7+ILYRaWAEDMxMogpmTOcAAsuk6HrBXHiBxjRAQzE8Hdb/s+ep+9DxuZwbLyfyIgIjKTiESEmcecTLSdNgAi0trGLMgcoxPxMjgLE5D3fnUtkenuYUYJIc4IZm6tRbhnlNIiwqetR0xEBpBEzJweYZYe7janyZqRtGnL/5IxRh+9r/p8gCCN2onaOaQ6izk5w1LdcRNqHEBYxN/85n/1Jz+ODg4ODg4ODg5+KTkC6IODg4ODg4O/OHz3u99t2F/v/d/4wWe/9+98onZiTSALx0PlIgPzsj9/GLfLnJOIMzDMVKXWwqCm5dw2KgVFs0rahFsCRAwCbjeKgDDmjDl63zOCiVqt5tb7LTM9YlpIKaxVtI5p+5geoaVspwYPJiqqICZm1aLKIozIzAg43G2O234dY9qcHlFUtloAynQPW9pZVXELj9i2E4tmgISJCEm0Jg5LXf5norv2FswZEb0jHBnpwQmmTE+bo++3ViqBrpcrWFjUA5Y5QSkagIe3Uotq3A9XZVEP33sXVVUtWhPkGW4JVdK6X/fbtV+u/XLr01Hbw8fny7/6w8/+2T//5++fnobHjz77/HK9ZuJ2Gx8+XH74w/d7t3wJf/HyPl4+Dqyhu68+9WWC/NNRMv3x17j0U1+UP+v7Xr70J/7vZ75cTgD01bfnV7n2nxV6ecOXN/3Hr2sSRKhUMk/3TF/VcgiWYeWrNwGEIIxSoAXMOJ+3169fnc5ba7VUfTi1T9+++Te/8RucMfr11cP57evHT98+VqGt6MOpCgHu/XY91fL64Tx7B7LWygQPu1wu2+l0Op8jvPex9/H6zSdtO8XL0iAxq7CoEMDCRZWY12FK94wg0Uyke84OBBUZt6vPKSqUlB5zzHTPyP12m2Pmqpkjp9mKf299T0BrISIWYS2eDJbTdpZSWMQjVcu2nbSoqggLEWWmzS7MtbbMsDn221VUSi1cKwmDgFWEvlzn6Aycz6dp081qbeFhc7JIWPS9u3tGMGgJpJHL1QJ3A5KZ55xjzjGnhxPQto1FAeruFpmEcn5sD2+3129RTj340vcxwxC7TVj84Qe/jfz+F3HooQ8ODg4ODg7+wnAE0AcHBwcHBwe/9OS3v/3Zp6ep5eOrh6c4vcGHUkrlcqq0NWXrMZ7Srvvt6Xb5YONWhB8fH4ULiVKtpMoicOcgBhGRZd58uFn4TJsCCFGGEyDMFJHhZhMRDKhqZpjPTI9EJElZVtjqmRHQ2qQUVgERMtk8lyzCggjCyIg5+r5fc3Wll306co4hzLUU/moqUESkFF2VVK6NmHMZM9b3ZLrnnCs3ByhzmScyw8NnTzdECAtlpDsRwq333kpj4jHmmjvMZNLCtep2IlWPEGIV4SUNYeFSPHL0voret733Md2TWf7wjz77F9///cv19sUXH3/4B3/0+z/87IsP1wT3Edc+n677NIvEZc4ZQYmIcPflpwYo15rhCvjW/Yu7LCN+PDP+8YbzT2bJ9DNCY/pjr3vvveU//dXw3Rb80xf108l1/glZ9r/uZ1PedSBfEgDoq2g7c5XpVVY1GGtEMu+K7/v7FUYnKEEEJvASbzOLylJhJJEyN9VXW1OA4KcmX//08Td+/dMmfKr6eDp9/dN3b1+98rF/+u7NN37tV988PqpQ7/201aJibiKkIokcc+x7P50ey7ZRrWkzzVdhmZAgyvAw01Iic792d8sIgOYcve9ugylL0efnpzF6LWXNZYYFEykrE9yj77uo1Fq381mLspLNCYaU4h4senp4xOmMUtmSWEg1phGRlLoa2Ywk4sy8PT+ZTSDdzObso4NfNCjMxIDH7H2/XlReTuYwE8HMiFhZMhHuPkxVkbnvXUWKqIebmZudH86qJcIj1+9CBAuXUk7nk6hmJAvAlASQEGtKST2hnmnbbn188eHps+fbrQeQ/+Cfzd/8VT6fqTf/5je/9Wd/aB0cHBwcHBwc/PniCKAPDg4ODg4OfonJ/NbnP/yr9KPTu3+C/+vf/rTMIpWqStuKhpMNshvHzjGIfPTrfrtkeiny8HBm8EuQGm6OuFcZmcUyr3338MxQonTP8FrrKkoScr2EEhATEROrUNW0mZlgJhZm5tX9BAkx8RIGUEbEGKsr3ccAkpki3Oecc0QkMdetZVJkIlNVaym8ltPoLoW4p1iAAxHp4RkZEememeExxiRmVlmCgntAmplIm8PdttbWet66smAWViYOEJhBvBbbmIVrSRaPVKkM3vd5ue3XvafodN9v47P37z//4sMX7z/0Ps3DPX/02Re//4N/1cd8vlzff/Hxjz7/+PS8R8ITHohcRxpOCAB5D1IBgJBJL2EuvSia8aUu46vo98dfw/7xHJl++g9+5oveZVD503mJeX+yovxnCKD/lGCaXkrMP3Vj8r6S+OWlMRNzLsNJxrorv4zGvwyg6adq4T9+OeuWJAgo/PKB4NVj+/STV5WpqZxqeff69auHs7m9e/34a7/yydc+eduKjH77la99+u7t61ZVharw4+NDa60UzXBmKafmo8eYTMjw9BkePsccXUQC6GOa+VJquPucY3X5S9E5Z2aUUpCIAJJEpKjWUpnIzJi51Lo9PKgKMTImKFk4zAGqpWatyTyvnYhI1GfPSBJ1s3DP8HU2ot9uZjN82VzCwqeHvbg7RETo7gxX1czsfWdmFp7ThEVLCfPMZFAtlZmm2bKsezgyATqfziIy5xQRFo6I9cO300lUEhmzI335QzJgkd1jeGZpru06vVterr3PGI4w/fi6t84BzBZHDH1wcHBwcHDwS80RQB8cHBwcHBz8UvJP/+l/S0O208df/6v/6Hf/t/9AyUnUMx6bPhY+adrlw7h+vDw9CVOrejqfhDNjklCuZNgNEQD158v+fGGWZE5ibVsS3fpIgEVOp9Occ9/312/eAPl8uSCTmUspRYqwZIaeT+XNqxw7IiCCTIRjDgAJ+G2HGyPT127fyIyI/4e9d/mRLLvv/H6vc+69EfmqdzebpCRapGUIXhvwTgvDgAHD8MKGtwMvZmUvDHjPrQ0DXnjlf2G2AxjeGL0ZG7JALz3SaDSkSDb7VVVdlZkRce855/fw4tzIqm5SL3ooUcD9dANVmRmP+zgRyPreb3x+XlsBBET0MEAkFg8Aljzsmpp6TOOYh5xSIklICOGhGqqmjcARos1LK6W2Zlp7DbPHbR4uIpJSU/NAROqKac5pKUtrbbffS05ERMx5Gqerq3APIMoTEAYgErmal1rDmodqDGnvxp99/vLTz7/44tVrDViq3Z/q//un/+rHf/nTl69eNQvVOByOy2JF18y4W4/jbNJYZ/cBeKwxqwdQ/8savr47xfhLVeMHRcU3vvuNevM3Pcp/Rc4cv9oC/TUQEYDofMP4psnjb3wo/2seuwfI+M3w/J12OXqojAhI754ifE2n+53fT/BhHc7XnxgBCMEDAEH4fEYY3EH13bMKgAAwQO/Z14ApwfWIj24uxkHI7fe/9zvf+ehbj68uxiz7MX/04Qff+uDFixdPDrdvXOs0Zm81tFGEa7W6WK1Wi9YaAEHoTE3NPVJKyAyIEQ6I/cWVc2biAA4gJOm+9XFcBymuAxtTRvAIhVAAAwhQi9a8VjNrrc3HE0KIcCvFzBHxPI3T3i05dzfrnnJAOlUtaoAkKaWUhpzHcZx2O2Ju2u7v7wEAiaGPI2TuL65hGKQ7Z3Iyc23r4M1hGBjZzWtr0zDkJP1jEmEuQ0YmIDi9fa1lTkm4v0jN7o+n27u7ubVq1tz3j55NV0+K58OpHdXAsXocr/SysDiK6x/9kx/+1ctpY2NjY2NjY+O3ly2A3tjY2NjY2PhHxk8+/thzixHiSumYPSIL3+x2iRisRpu9HK3cjVNmZmutx3Ds4dq0VSDwsGat1RLu45DLaSmnZZomJNaA6WJPzK0pi3DOMgzu7uay3wOR1gpmiEApISB6WK3EzEMup6OpIpOpuim6R3hEPFh6a6muxkSIgRjEqyuCmJAZkwQJcCLODhgefB6X11TdLSK01VZrqwuagbmWChDMhBDhbq5EJCw5JyJGImIiZAA0D2ROw2AIgcTDiCkhM6ohEqVsAQFEIofD8XCch3Gqtd7e3b56+/b1m7dfvbnzhvOp/eLTL7949fr1m9u5+FJjUb8/3B9Op+NcPMIDVNUt7Jy79p7ue+ksEkDv8faa8toTf7BtfD2A/qWo+b0b4Ln7/Es3+1W/4X4tOY51CuHfMoDGvymAxr97AP0uI8eva6a/liQ/fNEbzGs1um/FWhCnh9mFDzd9789+kBChO1cAkITcw9WBzr3zCFznZiIAWIRQDARDTkKIEJf73cU0jUky4cB0sR8fX++ePJ4oLAte7MZnjx8/fXRzfbm3tlgtHzx9vB9Hwn7UQyM8AhGHnHsWPI4DCyMC9SGPgIgCnJDFPVwVCVkkpRTu2nQpi7Zq1iC05+91WUyVEWutrRTTlpjHnN1VVavq+QhGuAMAi6Q1OU7MgiwaYIEe3arO4zgSrbVlQAwIQCJiFmERYo516Ci6OyCwSGvamiURZibiVluY0/kchbupWmuAaKZNa5kPpjUJCTERAYCbqzUP13BzwzQGD4oTDpeYpwZ+LNUaNsJBl0Bwt2j1P/qn/8Nfsag2NjY2NjY2Nn5L2QLojY2NjY2NjX809BmDyXQ4hV7OLMO4EwHGsH2C5I2tmS5tOdbT7XSxzym5Wv8wPqi1pq01SuIAzZqqQsRuHEzNm427CVkMcRwHZjZzTolTwvWz+eAigYBuXltEUBYMBHddag/5SimqGuFq5uG9ekmERExIRKi1gYeIEAMzCBNiAAQLI1EgAEkgeWAERkSomqqq1lrcnZlaa63VWgtGEGB0z2wft4YY4CwiKeVhQECAkCREBIHWBQIiwAKcgpMTaoRXc4MgOS5tKU3NXr56/erVV4B0P59ev3n7+cuvXn719qs3d63Ycqqvv3p7d388nE5LiWqhAYgYCOpnTQauleSvg2dtxBpAB3hPd2mVPv+KOBgf8tP+Ja4taUR8P0BGOCfRa/s7HgwcuJon+sjArzsq8N0zIp7T3DNx/v4akPr6dA6rlePr2/qutfxuQwIC4ry35yPyNYM1PmxkVz0DQED0PDogoKte4mFPEVc59Dk/h3eH+msP/HAi3h0ZQMLwCEBiiogw781zXNUs8HBcIwJhvfjRH6NfPpHznEMhmEa62PEgNGSZhvzi2dPnT55cXe7DWmj73e88f3JzNY3D5eV+HDMh5JyncdiNY2JixGkahNGtualb06ZIQiRO5GrWWhfHIBFEmOp8mmutZgoYiAGI2jQiRJJqs9YgIgsPIr027oQRCIBEFO4QIZJSSjmnlIREENCBArDL0xFRkkR46+4aIuLuh2YWBsBVvB0eHrVWMwNGt3CPJAmJwKGUYqr9dEcERFjT1pqptlZrrRHa/SrCLMyrrYeQGAHD3ALZgJYGkHcyXcn+2iWVaqUsbqqmdjoA8csTnhp9cuBtSuHGxsbGxsbGPxa2AHpjY2NjY2PjHwF/9i/+BbIZ04mma7hFNKTY79KTR3u26qe37Xig8MQCROAN6gnDQ1XneT6dllKAxIIUQPYXlAdHJEBhypKzcEqCIiAJUoIwXD/5TxABywwRQVDnY2hDgFqWcM+Jz9lumIUZILK6LaUEMxABYh7GPIwOgYhEnFgICSA4CwuCNwhDcCAMVS8LRphZqdW6NNeh1rqUYmYsvJtGD3czNZM0pGHk1B8Q0rngSTmjJGCCCABHRoAAD6jNaqtFATCQAngp9TjPVdFAgKdPv/zqi5dfvbm9/fyLL7pk4/Xb2zf3xzd39TirWdeWhJ/TtS6BcAQIjEA/t3i7WPlX/or5daNGIFK/PREAgPvXysKIiKu++ixLptUfLUyIABHm3bkNPUFlIgjQ8+MgQDdn94sBXUYRAHb2Lr/rUhM6QPhDw3gVfTAi9wl+Fu5u501cvRZn8YUH8Dnu7TMECTEiHIAEIcDNkQAAwh6eEnoA3U3c4fEu/EVERHdHBOyn8WzV+NvwcJf1Gc/qE8T1+++gb56Sdw/yThz97jv0nq+6zznsB4AQmIiIjiJ+AAAgAElEQVT7dgMkgmdP5emj/aPHj37w+9/76MXzyzE9f3zz/PGj68v9xZinJJkCrLb5YFpaWU7HQ69gq+oqLYdoTeelUPczA6i5unMSSglFJGWWJJK5jz4MIAjECIC8my6f3JSqHpHzQN0sjuvVIMQId2vqZgCYhgEjwky1hTsisAhEtFqZmYkdYlnKMs9I/QjgvMy1tYAQSUkEAM/ptNdS7++PkiSlhIiq1qrWWlVVPcZxEGF1ExFCbtoAgIXzkJHA3VIegKRozM1qBA37PO3zdLEbBwy/ffP29nBaSvHAP/4s/+FOHwHyif9oi6E3NjY2NjY2fuvZAuiNjY2NjY2N32o+/dE/L84OqdWJciOJKeN+l0IX9CVhwzZ7nbUsEEBICOTarJwwHN2hDx2LkHGkPOIwUh4xDZEHRCQA1kYAjASI5qbaTBUimLgPLANTAACM1gpGJGHpxUxrbh7eP5WP7iB5IGZAhJSBOcw4D5yz1oYAwgIBHuFuQBDopi1c3dVaBXeBqLWYtvfiRlxjvQhmSjkRExJ6BHEiySgcQBGQhswihNh0za6j2wfc3T3MCUjNT/PigU39qze3b2/vbu8Pc7Hb++X1m9NnX7x59dX9odTjfDqdTodlnktdajtVbxprsApwjk0BztFlrFP5/oYA+v2oExGJqKfZ30hAcU223xWfH+q8a4S6jmGENf9EFGH3MPeI6LXVaZyYWc0udvtxHM2UmYSZmD2iqQ4pj+Own3YAYGZzWZh5GEYWBgAzR0JiTiLjMIjw6Tgj4jAOhGTupSwsgoitViRKkrKImy/LnMeRmT28mVk4i7i7qjKzuy9LiT5c0iMg3L3Uqq25We/OE3OrrdVSanVfW+Vq1mozs4AgJFUzs28Wn+FdNftcbD4fOIB3x/Trt/+lh/jmD9//EgF+6czSezn16kdhgmnEYUh5GJ7cXF/tdzvmx1fD46vxckofPnvy7Q+eX07pajdc70dBJ3AKA3dwd9Vw63F8uKtZEs45pWE01aoqwyjDSONAQMSCw4gR6B5qva/sbpw473fN3SMIqefXrdSmzdSYERHCTGt1UyJCAHBfliXMkXCdiyiSUiLips1UzRwgzLS1RogAaG59eKG7AyAhE1EEmFn3eEzTpGq1NmFGYgDKObMwYCAxBLbWVNXDiSjlNO5GZgYk82gRhkB5tICmPqYxkO/v7uda7o+HpdlSIkHKL9PphbZ91DFtUwo3NjY2NjY2fpvZAuiNjY2NjY2N31I+/vjjK2mTxE2qd5aHMac8EMMkfilm8xub32o5WS3WmppFAAAhcg+KEpEwETESklAeB5kmGSZABk6RcwS4KswzuEFAhFutrSzaFAFyHqq2puoRxEREtVUESCLTODFhKXP3WjATIEFgSklSkl6jJo5mJALMdZ4pQCR1o0bT2tzU1VzdzE21FowQYW013JiJmZkIEVPO4zhQACIQAefEwuEByEFsAeah5jKOJBLuy7y0UgN6rdNPx6XWZhYBNJf26u3tUtpxXj777ItXb25v746n0r56c/j0s1evvzreH0qNXmoF71MBAwzAVxtxj3zPxdczXy/nrraJX+Fufu9LImRid/NY3RaIQEirrWKdKojMTEiAwKsLgfszpD6fjlm1BeC0m4gZIlpriJiTXF1dJ8m11svLq91uMlcmEpEeH9dWd9O02+0udxeAoKp39/csst/tiDkCzJy7JYFlyEmYT6eZmXe7SSSZ2fF4zDkT0zzPwjwOY07J1E6n426/Z5Gm2lwtAonc3UxFkqqfTqd4D3Nb5rlpM9NaaoSLpLLMy7yUWs2s+4trrafTydwhAhFLqbXWXve2CFPtvWkPN3dTC4gINzVfbdEQ8Ev15787v+q6Ar0XY58F3fjuawwQgAywH+FihCnRRx88+953v329G589uvrWi8eXU77YDVf7KTMKwsCcmJiRsK8GS4Q5yTBNZta0SR5kGGkcvWog4jiAmrdmrRELpcG1OXgwtl6Qd2diQlyWpSxLKVWEiRDCXZurrpqTiGUpbg4ApRRA2O92khIRqWq3vkSEmrVWc87MbGZdrWOmiH15MrOIcGsKELvdTtVabbvdlCTjqvYgJIRAd6+11tpaaxCRhnRxedHHM6ppD/IpD6W24/HIKK3o29s7HkfMeal6f5xbo+AUrIfrXV4MActIWwy9sbGxsbGx8dvJFkBvbGxsbGxs/Nbx8//rnxXgxfPLdvHtaQbO0zBcXu2mSTAKLHdwuqWoVudyuF/mUylFTR0wUPKwkzSyDPvdPo8jDgnAABwpeic61MLM3euyaC3etP9C1D+ST8RuxiwXFxeB2NxLaykPeRwP98dSm0eklEWECJlZhJmRhIARTcEsPMwsPFKP0TzaMgOEsJh5bW1ZlrmVaopMiNSVDeGhZvv9PuccEETMTASQcsrjAO4QjtgHxwVoi0ALnEtdSlmWKsOIRGau5ki8v7wMlHnRn3/y8vZ+boZ394fPv3j553/xk89fvXr99u3dYTnOeqpuHmamTdXcLPA8Z++9uLKPWoT3fm/867LM+BVV2/VhHu6NgLTGlHF2WaAwhYe5IwARSqKL/cUwDkS8m6b9fn9xeRkRqu3Fixc31zfTNH7xxRdlKc+eP3/0+PFuvzudTmbGgFdXVyKylLqm4RiA4B7zPLfW3H0aB0aqtfWm8FIWDw+AWs0telkVEWuttRZ32+/3gNCa5h5KmopI9wszs7CER+9os0gAlFo5CTGfygyAqd8YwNR7pZ3W6Xt9siAiomoDAJHkahCeUuqzDd1tWcrxeGRmRDCz4/FUShnzEBGttfv7O23KInNZTvPpdDz1zT4cjqut+Fyk76k34jd////bDGP8lbzzWD84sB9+RkAE7gAO3cshCIIwpjTllIh2I11fyocvnn/0wfOPPnz29Oby2c3Vdz54/vzZk0c31wgGVqGdos6olYUAMAAwHImAuRwO1hoKh7mr1taYJeWhauv/L7U11bMwph9hLbXGKtqGLNLFNR5uZoCkaqXUcbcfxjHlFB4ewSkDgEMgEifJQw6AcHcPZhYS9+73eDilmJIQkamaNjebphEBtSmY94s5rTVtqq1pU2sa3bGCEBhN2/F4b+FIIEMKgKYx5DGAlqVqBBDLuKc0oYynas3BCBnp9lqmo4G6U/vP/uv/8dc7oRsbGxsbGxsbvyG2AHpjY2NjY2Pjt4gf/eh/HXyXPe2c7mAYiIc8jLshMRNY6EnLydsR65wo0JqWBcIRIUSCJDjxuGOZmIacsjA5uls1LdYKuJIbuoeptWatgXvPjXplGCVxHlopECEps0ggLq1xynmYLMAtzIwlETP1Xml4hCEFCXit4EaA2pqrUUCouVq49Wyq1mbuSKThDkCJmYVYWCSIDHDMWYR7Rti1vT0RpnBtrSxzacVMGRGAgYQle0AzR+Jmfjotd8fjcV6a+Zu3h89fvv3k0ze396UqHOfl7d39l69ev72/P5zmoq4OGufxdmdFwy9bGRC7NxdjFTn89U3avzbMPP/iyURJaDdOKWVAGMfx4uLi8aNHHlFLZaZxHPf73bSbmLm2JiLTOF7f3Lj7siw5pZxzzvn27q7UMk07ZkFENTVVNx/HEQDKUlprbs7CAeHWbSymqkNKETHPSy+lqjYzNw8A7kaHlBIAzPPsboCQRNy91drdvuYuzMyEqySa+0DLPm8yIqoqMQFR04ZEScQ9AICIobfIEXt0u46hI/QIdzczIRKWcRzPEmxQ1dZazrkXct0dApjZVFutqgoAKaXS6lJKKaXHoMuydMlDrTUiRKTWWkpZlmVt3rauqXg35fDvyjc80esKOH8XEQCoq0ZWhTQRQlAEBghDznBzeXlzffXo+vJqN97sp289vfrog6cffevFo8vd5S7tE+4SjQIYjhAIEWbhHuD1dNRaIKLbqM0diYmTuqmZWjMPM++iDCTWZgBIzOoWAMw8DjmnhAAe7h6AGAERMEy7nEcW7i9vCyDh/lZAzH1h9I8XEBIRdedGBxGYCM4DJbWWWktEuJmpgjmYh4fWZmbCDBFh/k7/TRDgalWtqWnT6gCANI77YdyP4+Tr3rkMu2F3ozw0p6XWY9NmURSUT9DYPdpS/sv/7n/+Nc7pxsbGxsbGxsZvgi2A3tjY2NjY2Pit4NMf/fOmUKDcyetrfYqRiHGX0m4chd3LYT7enY6HsiwRygijYGIggGkcxmmk/R4lASdIY6CEEaiFNq+ztrmVpS4nCGUCQcQwVUUPJp6GMZAcAIAwZxqnOp9araqehsxJalVkljQMFxdCDKog3J3QrS6tLqUWAGMMbRUgEidTNdVo1mq1piklJkbCZVkAab+/pCQkzGn9zD6xYEqREpiGWyCGO7gDgDYtSyGEVuvxcLi/v6+t5nECTMD58vKGJGvEUur94fTVm/svXr764tWrL16++suf/uLHP/309ZvlMGtV0AAHAAQHsB43ExKTh3e/Rvg3J92tIXj3LSN6RFdYr67hLuv4JddGxMO0t7Xq+z5IyMxJeBzS4+tHu90OEa+urp4+ffLRR99299M8C/Nuv390cyNJ1Oz29lbNmPjq6tLMj6fjmzdvSim9U6zuZSl3d/e9Ixweqi0A3KzVWkt185RTRHh4zgkAWqtMHBGlllXja+4e7jCOO0SuTUUkIuZllpRySmWeTdXdWRgC1FSYegDd/6ithTsGEFMAmLuFBwBy321szRAxpdQHOEZPN3v6j31iJanq6XQach6HIecMABHBvI73G4aBmc18HIecspv1HHkchpyHlFPfiYiYpmmapq4AV7Pj8ehmOefT6XQ4HG5vb0+n0zzPx+OxqSKAuYf7QxDdHwRWTcg7m/SvvPDwzSWAgOtoSogAEkZEU+vLoptS3IzOwxvpPN6QATLB1QjfenbzO9/+4Lvfev7R88fPHl1+8PT60eVEYYkgERAghIdV1/6/5sRZBBA90FcFdiACMQOCmaU8iKTjcSZJu/1ezZAo5TwkYSbX5hEB6O7MnNNALNRHTzIFwFwqi+Rh8HAPgEBmBoCe+wdEa61f2mi1TybkVou7D3moy3I83J/muV+fQAvwCHM3Q8D9btcvY/VnI2JmZKE0iGqdl/nu/t7dRVIep4vL6ydPnhKCar2/vyeSlKbqgHnP08Wbw/Lq9nSs1YNM4PT2dtiNwOLC//k/+eH/vzfmjY2NjY2NjY1/C2wB9MbGxsbGxsY/MD/5+GMlZbFxaKeCAT4KXO4HIWiHeytH04IAp2VeSpVxZBYmyonGIY3TIEzEhEyADIDg3kpdTouZhRuFQziCIzpCADhRdKWwFnOLlAY1r2oGEMSUEidBIg0YxzFL0lYJkYUxHNzAFcLDzFtza6baWnPXcJ+X2cxZxMwjkCV7hAcMw27a73b7C9WGgJIHTAxCfX4auiGEuVatGKatzvOxturuKU/uWNWaRs7T9aPHy1LNYdhdzsXuDsvdYX75+s2nn33xFz/+y5//4osvX90vpSy1LrUd5+U4L6W5Wni86y2vVmB4J3IOCIz+JUZ4b+hGBAIiEKx5KQJEICAEMRKhWfT+qTsEABFE9MwcxiHtd+M4jdM07nbTzc3N9fV11zHv9vvHjx8LszXLOQsLAKpqn7C3lDKf5lKqmSMCILbWDodD7+qmlFprp3kupXRnAhIhYQS2pqrGzLjmp4CIiflhIhwidGVKd+92qTcirkEwRI/azdwDAoiJAEDNRFiEW609XAYAd9dWiQkRIXp/1t0dACgA10I9OIRDT3W7AYO62dv6c2B/2kBaPRvMHBGtKSH2ZLuPkTyfjlWcnXKGCPfosyYjHBGZOaesZgAwDLkH1pIEEAOAe8Ua1xPfo2UzO51O7p5ESrdK1+bhqno4HMqytNpqrW7e79cHWr6/cB5K06tK5N0QSlh3L84974ei/TrGct2Oh3+JIABBMEAimHLajcN+zBdTut7Js5v9k5v99cXug2dPPnrx7IMXTy92YyIYBDOjEEg/XIStWWnNPSTRfsq91Cw5dam3qpNIGgaSRJJQGFqBVmkdZxm9Ao3mYQYQzGxhHkEsrbVlnk0tPAj7GbTuRfeIWmtKMk270+nUWu1eFAiYpt1pnu/vD2bGLMMwuJqruXlKKeecUjp//CKIiSUxIxIArDG1ezBxTqm1Fm6IkfJARMuytNq0WW1KkofdpVJ2Ekzj0tppWWbz1ryNmRcFRQn+T/7bH/5bf9/e2NjY2NjY2PjbswXQGxsbGxsbG/9gRPzw1c++U+6u26snJS1JIGVIYGxtGgTK/fLmNYEhI5JUixaQd5ecEhIJRmIahtRHr3WLRASANq21LsXcIqLXdwl7NdXdFSmIiDi5RjiJ5EC0AAsPJFxTKjEIYWFEb5UAGEHrbFrCFcxCW6sF3MO91goBSKhNA1EkgwhK4mEKIECUNIzTNE5TmJubqgETEFitoRVMiUC1zvPJrbmrmwICsuThAmQwFG1BPIy7i9u745vbw9u70+cv33z+5dtXbw+vXr/58uWrn33y6Zcvv7q9X9Y65zlo9l92K7zfWY1V4Rs9OYWHiLK7nM8/698+qxV6u9k9ksjFbmRJwzBeXOxSysRChLtpvLrc5SHnIeecL/b7/X6/3+1SypJkHMfwWJYa540rpS7LcprnWmtrWkpttTVtEGHutVazHqGjaiu1dl1BQM+VkfqFh6Aulu65LQIKC0C4h7sTATMFdPlKYxFmIkA/SyiIEJFaaxFAJLAOndOeVJsqIYoIBJibamNhJvIIbara1r53PGSsCIQB0FqLCCLMOROye6hqRBBzuHs4rQG0iwgirk1sf1AqBwC4u5sjobDknFW1aevy7J7w9v8igpByzr2QO4wDAKjbMIw9ee+F9JRS72631gB6KTtUdVmWfuFhnhdtVZsuSzFTBDR3My1laU3NrIfRvQIM65WLXzGXMuL9f2kEnNfUeVAhrjLmHpPDOuaSAgiia6PHBJdTvtwPV/vd88c3Hzx98q0PHl1fTmOipzdXj68vry8vbq4uLi/2Ofe9MG2NyHcDmzZzB0RiIaSmFoBAxJIoCSfxZY66xFmk4+5hhuauDcKJ0Nw8nCUvpZwOxzCHAAx0d0BgJoewcDdNKU+7SWvVdW4kIlFKQ2tWagXENAzjfu+1uZoDpHHMKZE7EKGwR/RPBmC4mS6lABCJZBmyJGGZ5/taZm212+fDo9VaS7E+IJGZ00hpxDQ2zsXi7rDcl6WpVafBcsvNEuhl2kYUbmxsbGxsbPxDsQXQGxsbGxsbG/8w/ORPPt49+uL57//Zv/o//8M0GAJOWS4Ebf7q9NVnCTy0lrk8enS5v9gDMcgAeQAZgRkQoVVoLbTVsmgrgL3ZCREGEAQY5+w1ehZLqNqqVmIABFMXGVIahIc8jWnI7g5EJAmJAsEhWm1WK6hyOIHNy0nb4lox3HpgFwEeZVlYZBx3KaWch2Gc0sUl73aQMiCt+VyPdLsv4vYWIcJtmU/WSrgOYza3w+lUysKE1zfXF5dX0/6S847HCxovwfBwmF++fvvTn3/2p3/+4z/+k//nT//8Jz/95MtjCXWA98TMPfRzJOiRXvg3zAlfG0EX2HXTsX4XiSjcPIyQeuu134UAgB4c0WvCeH19+dGHz6+urp48efLRRx9dX1/v93tm3u2m/X6KCDVrrdVSVTXcl3k+Ho9fvX1zOs2laC1F1SICkdyjtYZI3W/QK+YAgIgsIiLE3NUQXZWAxAHobu6BQIiEyIFrHznOQuXeI26tESERaMcs50yIrtbz5z5AsOe/iCicHEJNSyk9FTWzHkAjYoSrWc4pJXGPPvEviRBSvPNrQO/Rz/Ps7kS42+0AsJTamgLAOSbWXk0GgJQyEZl3abh3X0k/3qZWa805S5I+TM/MuoC4az08fFmWrhMBAG1qZuM4qulpmXPORGymPfvuxVsifuDi4oKZ53lOKQ1D7lIYRlrKYmY9ni6l3N3dHQ6H0+nUt2cpC8Bad16X96q2frfCcI2dAxEgwB+uZXTr8RpFf93hEUHnax4Pdo4EwABCcH0BFxNNmX/vd777e9/59u9859vf//3f+53vfvvyYj+NYxJZjvfeFoqqda7LfDidLi4uLy+v5rnUWptpt5oMYwZT11JLcbNwW5YlzNaieHiE9ZeVR7SmrSkhYYBbJJGUUs7Jwrpjup+InFiYEWkYRpFkHsypd5Z5HOViD0sBd8gJUgIkOB6BCcZhfUVFWKnL6fTV3S0RD8N4MV0kTgiwnO60FQAHIGYeU4Zw0wbgtdZlWfYXl8jpMJdTaacW1bkRL9UOpVYLUFi+NY2vNJ1oPNAf/fCHv9479sbGxsbGxsbGr80WQG9sbGxsbGz8ffOv//h/E8pIFI4OLTHu90NosXKUqOSN3FJOyOjhOYsQwDIDADADoJu5NlAHc4iopag2JATC6OmRuZmL5EBa1JCEJUE3IAgTBhESM4kgMUX0/EhLCTNEVG0RAUjWqrYa2hCDAJey1NbMVCSxCEvuhmOWJMPAw0gEREhIBBHhqq0PvTNTNzPzWpu7I5GrQUDKAgjuZhGUUp4GzCOnMcnIMqjCZ5+/+vL17cuvbj/79OWnn7/87IuXL98cXr65f/nq9d394TQvVcHhbN0958Jnx0EfhObfMPd+TdwcDxaOtUULXaELAdDT9ZimIefERPvLi2fPnn7/+z9IKdVaaq0XFxcffPDCzCBARMyt94vN1d1arRHAIrW0WmsrFQAQydxqraVU6mqIdYMx1jbyWuxFIDPz89mBripGQEQmQqQAsPAIYGIiRqSzLCJMVc3c1nDQPZiJmWotawgriRDNrB+Qh9GKa/wYq/0aCU1VtRExwtmKHBEQwkxEZt5atabDOArLeoTPLd+AVc8R792zR/6rzgLfCZaFufscmJgRzbxfH2DmADDVs5oZ1rJ1ACIgEkAAYh+lGB7M7B7utmbBhH32YsQ50GfuOX4XD4sIAkZEz1J7yM5EjOxuAEDM5/GN1k0tiFRqOR1P/ZqPhx2Px9Mym2m3n59X37oQ3+k23mtGx7uc+t2K7EVuXG8fCBEABCDnznQSSIxCeHWxv9rtLve7Z0+vXzy7efr40Ytnj188e/z0+vIiY/YyJsTQ4/EoksZhZGJzrbUsy+LuOYswIYY2VdO+VJiJiVQVEFJK7uEQIhmIAjDnzMTh/WoFEaGIJBFiCvcwk8RMBB4sgkR9N+nsT29hoepmFmHhEJGJEdEimjY3Cwf3MLdiKpKEpcyLm2EAYKTM+2nU2lpZyrK0Wsx0nCYRCUDzMAcLrGZV3QJluMi7iwZ4quWo3oKN081nstyETvif/tMf/jpv3BsbGxsbGxsbvy5bAL2xsbGxsbHx98ePfvSjCYuEkh7HdMEpmCAx7pK3ct+WA4ILUWaRYUCmwAhw0Erz0bW6G3h4q60U6naNCFV1DxJGZmB0CPMw9ZTH4FQcSDKlhMwppZwShiMCEkCf7uYaZqamy+KthfXk1JnYtLk298bMklIz0wALTMMow5THCREJcRwnSNmZw81N3ZSsRVvm08FVw9Vaba3W2tScRKb9DoOYZNzvAqCZWSAPedzvG+elwf19PRzqmzf3/+bHP/3kk88//ezLn33y+edfvHz1+s19saJxzgHB1j7pGue98208JMu/bOD4lQF0BAJ2S/Ll5cXlxb6P+APAy+uLcRwI6fLq8vnz59///vcJ8XA89E7uzfXN7d3d6XRqTZdlnuellFJrqaUsdQHAIY+ttVZbK01SyjkTs5mWWvtUvYdRfITk4W4O0IUgbKa9khwBEW7uuI70Wzfbe/aK65i+1Uhx7gib2cPwQ0kizLWW7k/oto7w6DoRAPAIjyBmADB1RCCilFNrtbWWUoKAHl4DADE9hLauHu4pDT2Sxr59RH0DkggAuHspJSIkpV5SrrX2xWP+Lhd292VZkogQ9+oxANB5l0stqkrYH57OZxPNDRGFpdZqZj1B7k+KRCS8LIuZ4RlC7IIRd0cAYtbWVlP2+dgSIPW/EIlIV2kzc3eqIFFrbV4WwvWixf3h/jifIrzV0koxN3e3fiFIrR+3iCB4l0GfM/p1P84OcnxvXQaA95VO4ADgsF5u6a9dBiSIaeTLXX50c/3Bs0cfvnj60dPHTy7yJdcPnl7fXO6YkImFeb+bENG0HY8H05YSixATdmFLBOScWZiQmikiDeNgHgGYhwmZ4zwEsn/IwiPCQ1iyCBG5qdWKTAgQZl3qwsQYHt6vPJVlmREx3NU03BAgpeTm2pq25haAFADALOMowu5++9VXdakIQJnHcbi82FstdZ7n47GURU3H3ZTzKCktpaoFsQSAe5g5MaeUZbqA8bIRH4ovgebowKgVm0mz//i//59+3TfyjY2NjY2NjY2/G1sAvbGxsbGxsfH3wccff3w9IhM13j3h+wAZR3q0m9hmbgeoBxgEhgTh0BSrAqG7t1ZCG7oJWp1Py3xiBFPXplkyApoZIhGL9OGBwr52RBmRMQ98cQmckHitZHqAWaullBNAEIIQaqutFDPV2rRUCEcE6TIKt4CYpnG/v6BhwDzEMGIekRMEYmvQFBGaWqlNtZVSluU0jYnA7+7eMkISCq1lWeZlycM4Trtxt9/tL8dxjyKnpZzmMl1cBtGp6iefv/7xzz77l3/2l3/xk09+9vPPX7/66nC/zIvVXmI1qwAagN14/RAgByATvD8X7iGI/lsH0ASYklxc7P/gD/7dH/zgByllZiKCy+vrPGSzdUre4f7w9vbt3d0dALiZqn715u2ylGHI0LUnPU6GrhgOFjZ19zVj7ZoLNW2mOWVELLW6GQCmlBEJzglfv8/DpvacsJsjejgbCMSMiOHQe8YA0BNgOLeVe/SZc045iXAv5xKTqoYHATIzEQZ2m/cqYu7N6H7L3v3NKQGAqva9SCn1ure7ExISunr3h0iHeVmWprqbJhFBolIKAOSciWyJm3gAACAASURBVFYrSN+rpgoAIpJScveyLITERMQE3VmuyszjOM7zbGb9Zg+b2o+2mT0YmfujdbeGuTdttVaPkHMUHu7DOI7jWJZFVR8ScHxXSQZfZ/GtAXStVU0RMaecUlLTPudRRHLO0ziqa0CM49ham+e5lHle5nme6zLPp9Ph/r7Lo+nhesnD+jwvVQQ8p89wXtQREIJMgB7qED2Q7jdILLROwAyEYKJRaBROSDcjfngd//4ffO/f+8G/873f+91xGJLQxW4ah5yE59MpXMfEYQ3DcuKUhEXW2ZVAjuteAyIgcxrMo6kSEyD0qY8eoc20NTcXIjdrpfbif3gs8+Jmu90OCdx0nudSSmttGDIzmdk4DDmlZSm1lFZrX4ciOQAk58vHjwOiLMvdmzdaKwI6AjKmxAIggISg1qo280AkZolVfkJJmJFUWy2l1ra/vII0FCe6fBrD/r7U09Jas/FY6xDPfv9PLx6/+sP/4E9w+xfhxsbGxsbGxm+Y7deNjY2NjY2Njd8sEfHmkx+/vbv76Zdvv3tD5J4H2e3yQDBExfk2llPoCQSCoJQ5zMjBPFS11kqIhIDoZVlqbbvdniV5ELMwMzGzZOJEhJgTZolWwzTUSIRSommCALAId9WmrYW5Wx9XViN8HLK2NaRzczefxlGSQASnRMKAkXJO44ARAOEIqmbq4AFNQy0iamtLbYDkAM1sbWkiMJMwY3iftZaHKQ2jSCZK5nB7ONwflsNpKWpfvn7zk5//4t/89POf/+LlFy/fvn5zd3t7WJalqZudxblrCfRsyuhD6s7Oil5r7UVgWiOlCP/aGMKH6jQi7qbd9fXV8+cvHj16dHF52fvDOaebm5urq6s+le50OqacAqCWKiIRcXt7+/bt28PhsL/YC4u7zUvVpgDQDSe9/KtNRYSIkLCWau5JEp6LtxEBgEQYAee0F3v7+EF04d77yNFa68qDLln2cGEBhFXQgZjT0FqrtRJz33MEJERiKktR03EciQgQ1qPRD9Qq3Oi2lbU/vrqJ18Ma4YGIhIQI7hHhPZqUlFVVTcNjHWDngYhy1gEDgJv1Hn2vFff9dnNJiYjWgnNXYTCLSI+GPQLOno2+AWvBWZKbRgAzmXt4iHBEmBkRA4SaIawFXCRk4pQTAJppz7hTSnH2geScc8611taaqrJI72X3n66HxaPPKozzKYEAYiKiB3/IuY1NagoQ4zgBhJvG+aioNlN1VXc3s2Veequ91VZrrbXau/X5Ln3Gd192STlCdH30w0BMICKEszAlAgEIgQEoYBS4HODF00fPnzx69vjROMg40M3V7umjm2dPHz+6vHh8dfHker8TyOgE2s9Mt2ogIMlaRUci4kTMTbXWioQeptrcLQKYJRz6lZVeZO6HAyL6ymThZlZr7ToUYu6nrNY6DoNImudZW4vwJClJzimbeyDykNfrIv1Nqlb1rgPxacjTkHNK3fGu7t16QkwinIRFEhG5m9WqteU8BFJRj2Efw4UGza3d3t0ei89LKdD+i//mf/nf/9l/9Zc/+94Xx/zDzQ29sbGxsbGx8RtjC6A3NjY2NjY2foP85E8+np48e/G9P/zJ//1/xDgk4SQwMkxi0g5QDjEvXhZrC0DzqPN8BACm1FRVral3a0FgVDUDvLx6lMc9yRCIzDwMmdOAJOEGSSILlMXLYmVhYRR2RFQLVW9r5hXugMjMSy0eNg6jA6g59Al+SJcXFzlnc0/jwCk7ODABkS8nr4u3Uk4nrQXdvZk3h4hmVszzuOM8YEpz00DaXV/1EJaQUsrjOKiTmtdmh/vjmzd3P//F57eH+Ti3V29uf/KzT/7ln//rn/781es3h/C16fmQHL9rAgOu/ebVd+yx3uo8RhBpbbMiAISbIQARDUNOOUtKiYWZIuLq6urFi+ff+973Pvzww6ubmz6fz8NrqcuynE6nu7u7t2/f9rruPC/DkInoNJ+Ox1NZyvX11TAOhETE7tFH2OWcOUmp9XSa97tdz6y7+EJS6qkkBBCSkJi/s0z0VumqZ4h1dB0xO3hZSp+ZJ8xqpq3lIRNSHydIiPtpV2stpUhOgOjuBMhEKaV5nlXbOI49q+0P7B5dZMzMXdbBvGouuj6hh79+HnjYhRjuDhDU0+IeQKvCuX3c7/VQvnZ3JiTEB2tHj5iXuaS+nleNg+N5GmAtJQBSSqb64N/oWfl6lM4OjR7aMnNvoMtqHO5C5ljvizgMQw+Lu3+jV6fDHQCIuSuw++7LeZP6fZlX4XVPpc2didan+DoOYeaqTdUAICURJu4ZvYiIAAYT5d4rVzsej2oaEctpnk+n4/HYzNwt3M1M3fslFXxvPffXAQKeo+d3GfT6YnjvlufrPvEwvVAIhgTjSI8upw+ePfnuRx/+7kff+u6Hz7/97OZbj3aP94mitVparSklJgLwlJKqvn37BgBZhAjNrGkFCHdTrbVUANjtLwDZAxGoH3vm1K83ECEQOsBSW22ViPOQp90OANytlCoiTFRqiQAkypKyJJHcPxnQtKWcx2Ech8HN52XpInnTNg157FMiZa3J2//H3rv0SnZld37rtfc5EfeRNzNJZibJ4qNKVeoSLAnqbrsBzzwwDBhoNDzRB+hJzwzbaMMeamrAhm145oE/QHvkieFJQ7Aty265pFarWvUgS2TxkSQzmcy8j4g45+y911oerHMiL0tlSSWpYaN1/iwUbt4MRpxXxL387f/5LdUyFXAjAhFi5lDQgxo0dXdTb2bFtJo3A+rPqsFXN/ub62ls2kxbl/7oyenDfjDHp1O/Yug1a9asWbNmzb+KrAB6zZo1a9asWfOvJD/+3m8DAQNy85YgkWw6OemS2MGGSyt7nQ42jdTcap2mg0NFspyFWQBZW3MHYhFJnBIlAUkuiSlR7mFzAqpgSmaI7EjWWtOmpujuVq0VALCm0zSiO7qXqbhZkDVizn3HIkhopunkNJ2egiogAidevACqrbU6TlNQscP+RutErmCKZoxQxqmOlYkQCJjPLu5uTs9kezJWNZTNnQtiCcEvEgHSxx9/9umnn3/2+ZMPPvjwTz786OOPn1zejIfiY9PDNO2GYSqtVT3O5TsezFud0K/FX7I4RwCgRY7scOR1Oafttn/7rbfeeOON1x48vHtx0febw+GACCnlk5Ntbe3F1eXli8v9fm9m0YuNFwx4beattZwzM0/TxMwphXHYEHGz2bj79fV1SqnrOkpSSh2Gse+68BrHJEB3b03NVIJSArZwcwBEo7ksrHYBraBmBk5E4DOWjg6vmiKgiMSwwMQcO8spzc4KYo7Bkq3FBgSHnafhIdVaEWGz2QaEDbFG8OhAyerm4MwSBWCzcES7uyNxyl0887FFvcwznJvU7i7MTDCPnURMc/HZtbXQhdjCkaMYrq0R82azmaapluIATMQigbOPz89EQcODaIfnOkrWtdb4fjwg5wwAgZgRMQeABhDmuAcAYF6vCBoeZg8EyDmbe6sViXzh19Hh/dnrL9rJS3NcVQmBCUOHEhtMhJkl+uMi0vV933euOk3Tfr9XbaWUYRhubnaHw95M5xZ41NgJYyxlyJrtTyPweeQj4a1Rm9GGdnd0JwJhYAJE3oicdfkk53vnmzdfPfn1X377b737xqt3ToQR3RKzaSvT0AmD2zAOtRQ3lU6SiDDXWhA8JR7G0R3vnF+UqlOtwYpzzrUqAIgkQCShfrMhZiBUdWZOXQ7XByC6mZsRALAgMcSkQUA1VddlVSmuSWHJwOQO3mor0zSOu8Ou1UoAFxcXm81GhG+uL3c314f9LvYdF4uNVnN3IFC3ZlqaomSSjVKHmIHlMJVRTd0no+9fXXxze7hL+vf/8X/1Z3+2r1mzZs2aNWvW/KJZAfSaNWvWrFmz5q85H/72b3uPnrCBQcLMaduLgGErWHZtuNbxhq25Nq21Tx0h1VbMlRj6kw2LALITAREzo0MUWkEEmCEUCki1TNAaA6iZmptqkFOSmCtn0RT2YGEOZsbEksSJiFAQWASZ1J2SkLCVioicUjmMrspEtZZaSlNVNzWvWlSbmzKhiHRdtmZmkHJHzETUbzY595y6hmycU96MY73e7Z8+u3z67MXTL7/68MNPHn/29Nnzyy+ePHn65bOvnt8MU6sKhmAAc7VzYXfwtV/U/lxNaxRmoct50/fbk5M7F3fO71wwk4jkLI8ePrxz50JEiBgchnGItq+7TWXa7Q/7wz4MCapmFmCUEOahdYBLT9ksRMzTNMXXOWUHDzAtIuoe3mQiBgBVTUmIZgTs7jknArTFs3zcejX1hT7HbMBSq4N3Xa+q2pqHWwSxTAUQc85Bf1up4WI5Yve5/j03qf3ILQNiB8gGQBGO7irE6xLGdeLuBks1O6TZIaWwAM1IMxeOJjWGNnoWUyyJEZlLpRqIOOwos8CBogRty77O0wiDlcdTxXGeAXRrLIKIphp7hTGH0D0AsYjUWh0g5zzPP0wJAOYGdGBlM48VhcDuy4TG48bHoUgpHZG6u8crIgAukw9fXpRM8RJHu7ebLraM+bQyUZdza01Nk0hKSURmoYm7qapqrVVNVVsp0zRN4zjVJU3VYxDlvHl/6n2wtP2/9r35XeSAQOGWdmCABCAAfebzk/TOo1e/8dr9u2eb85N8ftJdnJ2c9KkXOD/ZbruUCFudWitAnlLqUkeIkqTr8jRVQDw9PVO1Uus83bTL5ggOjBjmEGLiJCx8SycCRCTRu29NWCQlYpmGoZZi2hxjGGYrpbTWUkoiWSTXOAuqrZRaa201/OMppc1mc3q6HYf9fre7ub5y05dmeAe3+R3h6MsnDAGiY87dSX96R5FL85txaE7NwSYyx6as4+Y31yr0mjVr1qxZs+avLyuAXrNmzZo1a9b8tcX/yT95ce9kyLmo2AVxl9S1I7yzAaoH3V9fXT4bbnZtqqfbLhFZ09PzO92mn8eLEea+JxEnws0GRcDdywSlQvBKBLDmdfRhGIaDaetyrrXUVg2wFC1VOSXJwikBsUju+hMHMI85bzl1HXTZXWE8gJkTQkptPNT9rowTIeQku+sbra1LKagZizTzpsZdMoCpFO5y1/fb0zORxJLT6QkxgxuoQjNrrqk3EJ3s6ZfPf/rJZ3/4x+/90R+/9y9/8N4XXzy7vNkXBQC4PVHtKL41P4I2AICfBX5fc3HMpDVkx0SEzER05+zs/r27Dx48ePvdd956+21miVl8XZenafr8s8+/ev785nqngTlVp2kChG6ziR5uKWVRSZCpxay8EB9H9Th4pd6aUGdqAMAS8wB9KBMAMks8v5odB9zFfnVdcrNWaozRAwibsyFTmKxD44yIpUwAuN1uQ/GMiJKEk0zT5A45JWI21d3NTphTkmkqRJhz1mX3mBkAa63zWDmAGIGYJAFArXVpZ8+9W2YGh1prUE1Ti7o3EYWuWlXN3BZtyBFeLyboeaAfEWlrbm15GCxMOZrEnNJsxG5NiTgv3e1SioiwCNwaDBgAuu97RBzGMahx0H9CnKYJELucVTXMG7GdoX+BuZg8KzhssZCEe/pIzyGcHu7uPutIQoriPlPvoxjleCkiIpO5x5jEYNDaWquN5ydAc2emvu9qrbWW2Bitzc0lpZPt9ugnOT072W43h8Nht9tdX18fDof9fr/b7QLFHjfc/ecA6J/9DxoPQB/tbAMHdGcCxNnLgQCqwAAJIRO8enf7xmvn33j0ypuv3Xv91TuPXrn72r2LV+6cEoStemLmnLuT/qTv+7i6ADB3HRI62FSmwPrS9USEtYarYxwHJJSUOIurtnEsZTLVtIhfhCWnJCI3NzfjOLRWAMnBWyvDOJRS+r5nFnccx7HWFkZyZtlsNkjU1G5urpn5zsW5MJm23W6n2tzjIiQijjUDN4vFPElJzdSMMJQ2ApQonyDnQ4Wr4TA0r+bT5V3Z3nBu/+A/+m//gp/8a9asWbNmzZo1f3ZWAL1mzZo1a9as+evJ+3/wv53tpwefv/jg2w9cKCc56ZNApXaj4zXUAVWZxc1dTQjRAcwlC6XkzEAUHUtVa2pGaO6qzat6UzAFd3cr04CuiaDVAm7CBOYIICkhMSATM/UdbrdBcxnQWYAYPYgeqamZgrZxHEqryBgTD02bm4IamIF72HwRMeVESUiEut4RWm3c95Q7YjFHc3RiBwTwxFJLvbncffLZk8efPf3iybP3f/Lpex88fnK1u9ztbnb7w2GaagvKDACE7BAD0OZfyfwlfAb4+QD6pY8DARDp7PTslVdeefT6o4cPH7z24LUuZ2F2cDOrrV1d3+x2+/1+L8JmNgxDa2oGzKRNSy0xIRAIg8+WUoJvllIJOUbVAUDXdWpqauZGRExsZr4UXWPq3UxULUrUICIUEHORbsdougCECMBzKRgsZqzFJEA4ukM8AKyZB7c1M8e58Orupha6W60BQKk1BQSOmnwcQCIAjF2IjvPxH7hV3Z0FF4TLvximFlgU1XjEzWYejfsQkgQbjS4qALwUZTBba6rta+duPgjRsY4Rf1SmYg60zJAM1uwAcTrcPYYHBn+fqe5Cun3xTSOiMMfWzscZ4DhX8OiA9oXjHvdw0YdjHHE1c7PjwoCZ4bL28DPTLJcLlI7rJUTxEm7RVYfZ70FELGxqZhbDHmPCIRElkZngE8zN6JcXOcbVMozjfr978eKy1tKajuOoX+/O/zwA7eC++KHRzcE9avxx7YRo+iiM3iQ+7dJZn++e5Htn6e3X77/75oNfeucbb7/5+qPX7nddQnDThu6gbqqtlFZrUwNyRHDE1lqtFQiZKBETobZ22O+QcF69MNNah8O+lgIAm82m7zt3qKWWWphZhEWoNW2tNq20mMFba+M4IZCI5C7HNUlIm82m3/TTOJVSaqvb7abrcrzHzeJiZmKJ9RwmRiFkCqeKq3qsw7RGnADFII2Gh6JDrZe74aY1BGZDNBKnf+8//S//1OfQmjVr1qxZs2bNL5YVQK9Zs2bNmjVr/qp5//3/maq4ildJSWQriUVQN1iT7aHty7j3WtCs6zahgHBVcCcEADW3aqaOgMhRvG06kz41VQMHmm/299YqBdZBDOEsARCSdGkufDJhTtB3UBu06lUd0ZCiqOuOtZR5ElqZmjZiCmWwm1lr1rTLWUQCyxGhJObEzByNbKsNJBtxbQaUDGWsehjK7jBcXl1/9dWLp0+effTTx588/uLJl88//vTp4yfPRwdDREINPwFggFtCDgnGSwDtftQ64/L/t4esCXO/2dy7e3e72Wy6bntycnp6dnZ2dv/+vbt3L87OzmqtwzDsdrvD4XA4HK5udgGgiQjATY0lhYhDVVutM1SGWUYcZWFCKqUyS9/3U5ncXETCK6umzJwkNW3gRxo+z98DACCsrdWqOadZ3wxzczNawqqNEF/Cx9BlwGL4DURpHjpjAGgtespsHoZgi9mGtdYQYNDLrjAeTRrxx2MFOHC2uyGRsBxZaux1ay30CDFMj3nel59xGc+yZrXSNOd8tC27e9d18ybhbLZwMzeF2fVsiDFukGptga1FhJlLqUFjo24M7uFAEeaAsMJs7nMVHVFEoj87XzBLKxgRA5jjzFkRogBs1rQBoMT9BAv/hoU7W4B+gGjKH2F6EGckig14uTKyTEeERRrjbu4Q3XObZSk49+iPehOYXyv2YrmwcR7tyLPnZX4zMseoRgA0t1rKzc1NbVVVx3EML0er9Tj88NayDILb7J6YLw4MdzfM60+wCKbh+I7jGFcI0DOcZHhw/+z11+59442Hb7/x+luvP3j9tTtn29wnTODsTu51HOo0RvEZmSRnVZ1KAfDA4cIMCMGaiVCbEpIkqaVoa47e95suZ3Ofxmkcx8120/dd13Wt1daaass5d12OK7NMU85d7nLuunhfuFnfd5u+06ZlmoZx6PpI52b60liCqoaxmMHuUcRvzVq11rS0WhsAmUEzG6s3ytKfXN4MX+0HIq4unbJKczQk//f/w//uF/upsGbNmjVr1qxZcysrgF6zZs2aNWvW/OXzye/+rrJabno6yLAxkpy70213sgWpexyvoRVwBXSvE9Riba5dmlYCEEHXqYz766vLUtQAN902BvepRYOZqjoQb8/OFEiBct+TJCDqcp8kiRCYITgkhlqgjCAIaOANavFSvNQa5UkzRwLkcaq1aXNDJhKRlLuuSym7zhXQ09PzvN1CyiGRRjKwBtpAG9TqUy3Np6rDVPvTC9mcXe+nz7588cEnn/8f/9f//cc/fO/x4y+urqbD2NTdwA3AEAzBfJHY3tYIhJYVGWLWHcT8sbngbACEwAQzWCTcbDYPHz7827/xG2+8/vqrr7zy5ptvAtDV1eXNzc2LFy+ePXv29OnTZ8+e7ff7lNLJyQmymHmtlQjdvNZYIkjhJgYAZiIiIApWG01bZkagIKmhA66lMjMSxtQ7Jlabe7VzuRUxIK/kpGYBsgNxhuYiHhDSCWHqco6heYTEwoBYW43iJiG5z8/wM7+sNm1VW1R0tc1YOUtSVTPNuWNmIoymb1BjIkKct2SaRgBYwLHPe7o0oImwlOpuiJSSIKLqS60zEREhADS1cSpRUaX5IFE857j4MWh+VcC5HluO3x7HsbVGxAGgzZxZksg0Ta01AEAiXArggBj0/HgYIYwlywBDZrYQjrgHnYeFqh//xVZb9NbjIIRbWVW7rmcmMzuKqltrqpZzcrNWW/Da6EEH479dgkbE8DmotsDNzByylNg7ESmlmCoBMAsATtNkNis+4NbwxtyleCELgXhrkhIAtNZOT09PT09zzsyE4GpWajmM4/X19f7m5rDfu8XAwvgfgTcwA7d4vzBRzFd0mx/1cranIzgAGi4TPwmAABhREAgxEd077X7ju4++89Zrbz26/9r5yb3T/s6ma9O+TUNtzRyQpd+eIJGaAmBrOoxjkhSTCdWsTPUwjF3X3b1/L8XCHFNrLc51OF26Luecc0oxa9PMRTglpjimxH3fifDsIAEncNcGWmNnArLHckuU65Gp1jqO4zgUVRNCg2I2aSu1jLVM1tQVXLHW1tSamxMZijrl7R3pt5VkrDYZujqJautrlTZ0qxh6zZo1a9asWfOXywqg16xZs2bNmjV/mXz427/demDCpLnkitm7rj8768ArlR3Y3sfBpsFbtVbdGiMyIr20LqhpNa21HLROMFcUOaeekBxQup6kA2RFAhbpOyAxEpaESA7EiKFfQDc3ra3U8aDTgOjBe9s0gLYsjAAO0NRCCo0kBtDMebPhvkNOjEgO4Og+SxgQCJnNzbypV9WitbapoGPmnPK2Kjy/vH52efPkq8sPP/niTz764k8+evr4ydOvLq/2+0Op3gwc0DAI8xE+L4aHpevrDtHNhKXK6nNHc+4+bzf9nTvn33jrrYcPH9y/d//s7HR7crLp+5gOB+673f758+clJjC2Nk2llNJqk5Ryl3VGsWA2exSCe861UMR5zN7CFueJfQ7ui8Fg9kLMTuFaKwsnSbXVYKBz5xfJAkeazhMLCbXpNI05d9FZDr52rM7SLKj1KGxabKO5iCCCqoYOehnuh0RUWyu1iAhx0F306CSbI0LOHQCotqDPKSVVDaAcjwwAnVJurbm7LC3suR5uVkoFmL8fT3KsDAdrdndzULvNYYkIF2HISys0uCN4lHxVw0YNHhx0tl/E43E5gOjutjzPcUjj7eGExyePLVkukpDVKGDs6JzWNKbhxbYdhw0iUoDM8FBb1ModmGk2PFDMwpt9HfFaL196uVZja8xj7+SlSttjNWIe+YjHq33WZLu5EZKDx3RERGRhM40/xitH+b3WOl+u7uGpmFEzkaq2VstU9vvDMIy11mmayjQFVw5yDgBM87LHPFbyeEMBAtjsAwEAxPnGBDjKbQAYYJP40d3to3ubR/c2r987e/3enYf37zy8f/Hq3fOLi/NmVmoFJE6cheOiIiRAJGKJTyokNY8GNCI7eG0tPOCSBADcLE5uKSU8JA5QpmmaJiQQkSSCcyN/fnOieytjGQetdb6BAZCIJSVVUzNA9NnTIuAArubFoaCrazWt6IjABAKA6la1UUqAOE01d5t+e155CyLN6PowjkUnsOGrs74fOtbVyLFmzZo1a9as+UtkBdBr1qxZs2bNml8s7v78s0/GqxflyfPxAnqClFMiSgm3yWy8bIfnddy3MmltruratLUkKeUcUCZuhm9ap/HQ6oQIm00vLITCLHG3ft6esGQABGYgcnBkAU4AqOqtKiFYa8NhRDdXnaZDLZO1CmCELohNC4Fvuo6TIHFMXUspS8pIrADU9ZizI4IaNPOZ5lEdR23qDg6mrlVHNVUzbehGDtKUrq4PH3362YcfP/7g48cffvTpTz999viLSwUIwzESA5IBBvjy2e3siLcZ9Aygb4FpICAmZOF+02+3m+2mv3v34tVXX33nnXcePnx49+Iid52ZXb54cX19c319fX11eX19vbvZmTsR5ZSJGJHcnUVYuJQC4NG0DSQVPVw4EtSgcIgzL5w3FtTmVuzMpc1j8UC1xfyypho4lRdtgrs31alOSCjChNRaPRwOKWUWMdMQ8xKRqWnVlFKUN2cHNKKaqs4OYjMlYgBvTcOPgUi1tdrqceRdvGiZJnBHpJxT1L2Dt95WZERCykzEsIz4i++LcIDmWhsApCS1zpaMxaEcV34cMYzL6chtETHc2V3XLd93nCn+nMC4rbWcExGrtvB7IM7Yt8uZiNpSW17ODLQwOIuEmgMA5t0HOPq13V1bIwmXzEwrVfVo5IiTHpVzkRQN7ZisOCuDca6Kx8kGdwK0Rd59ZN+0uE6OADps4yKJCI9nys3VrLU2mzQsFjY8jMwhg3ZwbRqFbxZRbdpayE/i6gUAbW0eZGl2BNCSU9d1KaVY87jZ7fa7fal12O/3u52GBERbK8VNj9Jn85enbwbMvpSgwec34Ncd1wQgABnhvIO74fThegAAIABJREFUW3ztzumDu+eP7l98661Hv/TOm9/+1jtdl5EcCXKiLpHWAu7CcjzjiIzIyBzuIDdvTacySUo5Z0lpXoswL7UcDoe+75Mkcx+GYRxHd4sSd9PqZrOtBgEdWpmmcahl0qZqCsTC0nVdbdZU46xJSozJ3bVV84rQiBxByT1LTpJFOiJS99JKyhkRh+GQOKXUD1PDtOnP7h8UL2/2L3ZDbTUrP3O6Uno69b+1VqHXrFmzZs2aNb9IVgC9Zs2aNWvWrPkF8sN/9s/u3L949K3v/OT3f5fEEuLJRs42jNNNPTwf9y/K4bpOA6FFHzYkBeDIIswJUdwREPP2xBwOwyF3Xdd3m82WJCPxEQ8hIqpCmQDdrfkwQNxsDjAM483NTdd14DAcJgNzB3MXEUkS7cKUJfediKADpgRJ3AG1QWsQXVGR1lqtrZQaZdQgfUziFhCrcSJknFp1Es6b7en9m4N++vjLP/z+e3/4Rz/4w3/x/WeXu/1Qa62lamkKixU3dAdRe7aj2BjA0eYCcDQxfZ6IhjD/Q4hdl+9enL/z7tvf+uY333rrGw8ePLhz587V1fWL5y+ePXt2eXW13+9rKe5gBqrtNmk1tTbDcmVmFg6nRDBicw/jcIyHmyvYZnEbvwgDwFQKIhKSmduiyyVEJLKFA8agMyKCWdEwCyI4ppzNp14JZ74ZTDaavDGVztS0tqCi4W1o2gyi/DsjSABHJPe5GcoiwdrUjIUBQNWSCCG22m5LjeGW2VlEkLDVFuy167KZT9N0cnLCzOM4RHW31gIAx0J01IcDTAe+JiIzLaUyMzEDzm1iZhZJzHRzc2NmYYIOli1MtDiO57PvbhazB2e5BxESpTBR5JSISM2maVLVvu9jiuM4TYiYU7r9NkREYo5OcSkltL8x8m+pWvsRhS8N7jiwgAhhdlC1qAkTcSDpQOGqDQEYiYgcwFSP/pCoJ0MISRDV57Z+PHmYWBDI3N3c3Pu+T0miFxxN7XgzMBMg2iL66Ddzoz/c6yHFDh5ea3X3zWYTuDws3pwkysLzMEx3SVKmKXTnV1eXz58/O+x3ZRxiQinifBJC17G8++D2zQY/79POEZwBMkFPkIg65o7p/ln37puv/b2/++u//J1333nr9VdeOe3YoO4ZVFsZh4MwJxFhKVMZhwGR4ny02pqq+1wYV1Vzc/OwsgBCThkAx3Hqui7nrpRpmqZxHKMOz8zERMRMcw29teoOQOSIzNJ3fVOrZki43ZxsT04Ph6FMU23VTQFNyN2diS7O72y3Jzl3bt5US6uShBDLOAESkxgwS055s59sX/T51c3z4TApqrfvX118Y3s4k/qb/8l//Vf9cbJmzZo1a9as+RuTFUCvWbNmzZo1a/5C+d73vtdBE3BQStK6vtt2Alao7WC6pLqHsq/TXmtx05SEhEGEUkYRIImxaGAIQIAkKTtRdWAiDqewgxkgoWprraAbubIpuoJWHQcwQ4Sw4tbaUk5E3NSAyJHAiUSYuZkDMSeZNbK1zuATgAEIYBoOCNBtOvcQCET3GczB5npmNHqFu+RMpdZnz68+//LFk2e7jz599v6ffP7x4yeffPbksy+eDFNR9QDHBGSuM7KNwuwRcC2Ey8EB/RbywiCCm35zcffiwYMHDx88vHtxJwltN5uuz2aWc+q6/sWLy+ur65ubm2EYQxYsKYlI4Dmce6no7q2pqoVkdymZzi1dM2+12qKLnU9IlFsJCQkAZg0xIgAGRrztODYzIgqyeXQKB0DHZQggJ1LTWuvig4DW1MxmkI2LBCGsDqEfmVvYELx0eWZcarMQW6utBR5WC2Uzz1Zm86PdGBHDPmymwzB2fZdTjql9ZhZAudba930Yn49uCoiBk5LcvZQSCDu47WzemJ0GAAA296dfPiDsyUfWjIjRgDZTRFoa1r6UqeM3cAeAlDpwaEtTG2/halpochg2cCHsR23IbEdRjTWPqCQHRo9ecyRk0MdmNCyzGo/t+NgXIopVDCIE9+NRnV0kce6Wenac7NlWsxxAZkYkAFTVOLMss5rD3RGQhcEhViPmLnzAcZ7VIUlSbDAARI8+rt6cs6rWNsumSQLC4jIQEUVETcN2Hesf+931eDi0qUzjOI1jmaa5XX77rfdycejWoM+XmTvSBMCzlAMFoEt492z7zpuPHr12/+Frd99+4/yNB+ePXjm7e77thbQVUEWwxKSl1mmCeRbkbJKJ5ZOow8fGHw6HuDjjFIzjmFLX911cYGo2m8znSwcRQJKknEkY5zseLAYiOnPctiCSRFKpRZsuem0DMDcjxL7rEVHNY3ziMAzx7G6xfOWAJJxTtxmLToaDQnU8qFYFIKhqGyJxoIarkWPNmjVr1qxZ8xfJCqDXrFmzZs2aNX9+fvJ7/2tBOWB3ByZJAEinfXeSpe2eTtdPD9dfJrJEzuhIyMw5d9J1nLOnBJKcE5qBKqgFgHYzZMGutzppqbW2WpuqMUut0zjs0DURdMJoDbRZK24G7kTMIpJSlECZBVgcGYDc0QCm2pyIu87UWmvTNLo2cJ+hNMt+vwOw7aYjEWQCQjdwQJas6lOpLDmlLnV9ARhb3d3sfvyTD//w+z/6/X/+gx+898kHP/2yARggzG5cQ8CELEjqLXDwsRkKAMd7/uMmfwd3BCZm4ZRTSrnruvPzO6+//ujdd9/95e985/69e8PhcHX14ssvn37w4QeHw4AI01RMLeBbENLcd13XHYahltJaE0mB/5qqm6WUzF1bg3nKn5iamkYvNQB0IKemGhg4NCFm8xREJnF3VWMmZklJmqqpEZHDsnMY/WiK/rY2NbfcJXOrtTk4Ih47qsx03H5CFOZoNLt7DGcDxKa11SZJiBgB1AwRcs5mFhQ74OM0joDY9/2ML2GeJTiOIyKmJMysqsMwdF2fc4Y48u7RawbwuaJufpRaBOwOh8bhcOi6TkRaq8yyuKQdEQNkq0NKKaQWAEBEIslUx2kZQohkpqYt5MUppSMsjk40EQfLzblDwNjapsrMXdcR0TgMDsDMXc5N9XA44FLwDqXIUlg2AIi3QtNm7su+mMM8R9JMLe47CMV4rJHMIxkxpRQteCZu2kwttlZbg7krj7FW4H5cXpl11UdwXGp1s67riAUAaqkOwMTRhI4gQtf17lZKrbWCQ/TTwaG2RojhFo8Kdpx6Eck5hau6lFJKiVmHwuzgptY0yu9ISwG87/uT09Pz8/PhsB8OhzKM+5vd7uZ6t7uptQYKn40g5v6yEX3MzwDol4sKAECADORgBJ4BGKDP/O4bJ7/y7Td+9Ve++c4br7567/y0z14n0Cpk84devJGaIrKk1PW9maupmcXnwDSO5iaJ3aw1q7UiURLZbDYpJUmSU55hfdyYYCbxwbHdxHRHN4t/F1NCEW+qqqYKi4AFAMysteZmYGZuwzjt94OaTtO43+/dDAGJWFtrtYIjS865b+ZFYTJIZ/fSZuMkxYpWcC8ykHNxa9Lav/uf//d/3T9z1qxZs2bNmjX/WmUF0GvWrFmzZs2aPysf/dH/HtPUWmnG1GXciHTsVA467tq40za4VUmcc+o2PXUdpERA6I6qbZy0NXVkJkLQVkOPa60QYc55GA/DeDgMI3PKebPdbN11mkYiS0x9l1wV3JBoRm15g8hoUMrkZsRc1Zo5GNZaS63Nvdtuz+/fn8ap1QJuSSinxP2WEFHNwEyb1dKgVVA1UwOgdH5+L3UnyBlAxrE9v7r+0ft/8sMfv//jH//kp5989vjzZ5fX+5vduBuKz1AKZ4Fz1D4hDANhdH7ZhCWIwXR4+/snJ6f37t176623vvWtb7799jspp2kcX7x4Eb3Iw2FfaymljOMYGM5sbqFGAXwchpRzznmaRrPAqeCAc63TrTUFM5j7qSQirbZw78YGhBWBmFXbPGsOZ7Tt4ESUJJtbrUVm20GapqlqyzkjYHDP8PwyxT8UUxBFhIURaRzHEHHknJlZtTEzs7TWCDGxhBbjODfv6OtIUV1vjZiQ5kbtUmEWSVJKQcDc5Si7BlV0j/KvRfmamaKZ63MbVBBxv9+7W0rpqA2ptapq18X0Qj12fgOXx9eImFIC8KXmjMwS7dTWGiJGT7m1VkrJXRaOGYYW8wwBYBFJY9ilY1pdSpIkEXEYt+NoxFNFZm4b5wt8qbFbbEbsICKGt1pEHAN1anhCVBsTpZTi8eY2I2xbtN6hFwGIs8/CcZyXuXxL63lpW5dSFhAf8waNWdyhlGKm4BAH3QHKVNyNmKN6q25hjmAW1VZKZWJ3iHPNwu5g2sw1/NTgUGoxUwBMSeLcxblQM3APm0e4To5LIbHAQ0icJOWu1eKqiNGTx7kFr1pKmaZpGMcyTVobLPu4gGaf71xYZofe/jCM2zcAHJdONBFuOz7fdvfOtt/55qu//K1Hv/JLb9+/sz3tJUHzWry1LiVCcoOpFAfabE8kJWGWFDXlmLJoM3YHSF2KsnuXOgRXU4oivCoBooM1jSW7GApJREJkquMwxijSI2BvTQlBUoptKLU21ZBk19bqUW5uFgCfCYVFeC5WA6Kq12aTetqcyuZUkVnYrN7s9oexFNVuGIdTLX218+E3f/N//Cv9sFmzZs2aNWvW/Osb+f96A9asWbNmzZo1/z+N+289e/zOdHiu4z136k83fScMim0v0x7rSFaIDVKH6ZSYmIlF1LFNqm3y2rxUrxXcWcSJALy2Cd0I3LSgq46o1shaJyaCOVEmMzNgcHd01QYeN84Tu4E7ujckZOSq6I4EcVM7AgMwQ84CkPs+iXjnRAhak7DkhMyqHiTO1FS9gTtT2myFklOqmHf76Xp/8+Tpi08ff/nhTz/9k59+/OFHnzx+/PnzF1c3+wGAzMFuHaHjVxa39COEOGI2UoR2Nu7zRyCii4uL+/fvv/baa3fuXJyfnZ+dnd6/f//87LxMU53KYbcfx2kqU6klbAxJcvBZZoIF1Jqa2Tw1UCRFwzFIYsikzc2hgBEiMkm4NViAovkLs3mDKNQnfFvpQEzxNTODQ04pCBcTW06oJCKI4E4xoS4eGSaMKOKGQ0MkIYKZHdvWRHMTWURi9trsgBY+ktZFfSKzTRjJHVRrPInP1g4XZgCE4zoA4uKOoPhj9JpDG6JqADF7MIQPxxryUQQy96CPkg0RqbW521E+YabzHDkP3/HMxJdX13hRd9emwcPNNJ4+nrmUQoQAnc4EsJrFgkXzxaoBR/vEYkcJHEyExLRARY/Decs+Qcdhgz5fhS9NJrYMC5xHXmIUmAEJo4Vt5ricR5iLzvN3jgg6WDwRqQb7nik5s5haqDmOqBqJskjUt8Fd3dpsOCGRpNpSqil1CNh09oADoFkz02DN7p5yMtPWWmxYNNzj+Jj5ct6iCU4LQV5GHRKhAxOHGkdEEgshOoCb1VpLKVOZyjiVaQrjdlg7fFasBH3++kTC5S8MZk3K/NfmdWi7oX354nA9jk+e7z/5fPfg3ubBve3rr9x59e6d+3dePTs5ESJTK7U6QEpZmImREFmIhRDJ3AzJazP0WMBQtTZNYG6mYTsxVXQgBEFqtZWptlrVzMGi4Xy8aGGZEtlqDZdL67qwqMeFQkRdzj2iJIlNIUBEMFNCFGJeXChqpurNHRgBRjUU6PKm2xBe0dXVvo4dayV77Vqebv6n/+If/oP/7H/4i/+IWbNmzZo1a9b8zcnagF6zZs2aNWvW/Jz8+Hf/6dn9Lx9950c//r1/hxNt+v70JJ/2bLtndfeVTwdh7HIGYkjZux7cvFUbp8PusN/vyzS20rxpStJ1/fb0xMG1tVJHQk8MYM20aCubbe76LnUdcucg0FRba61EY9Hdwo4L4GqgBuYxbWsLEHZg3Gz6rssAAClB10GIas3AQbXVYYimojpPpY1TqXVycBYCxrzp773ygLttNfzy6fOPP/78vZ989Hvf+/4//xc//Jc//GCszRGFxdzULLEAeGnteNO+48tfpY4lzRmBEaK/1PWGh+Fvfee7v/arv/Z3/u7fubhz4W6fPn784qvn11dXz796PgyDuUV39dhTDvlDKRUZYRH1gsNUplqLmYYIYnYTIx7tyrVVN0fELNnNS51HCxITLFuFiEjoSws2SLcvRun4golrq6YG4Wh2d5/RcNgnRISZEaG1FphymkZEyjmLCBGa+TgOqtp1fWu1tZZzB+6tVERk4ZxzrbXVBgDEJDxXhmutQKhmpUw5Z5FUygTztEMOgYYvlfO4WuJvRSTsxinlmeECECEAtlaPqBdg5qrHnq+7h0U6pVRrdEk1FBCt6TyXkolZcu7DxB12iChBHwlpvIRqM9OlHY7jOLpDzpmZzGwcxxhgaOoBBKMrXWuNQzpjcjOmWXYdvWkACMdIay1oOHMA3JfTLltrZhbukabtiFLnqxHiBen4zVkaMnfY9bgvy6VLAakXoK9xkEUEkbTpOE1HP3WcHfP58cHlS6ux8V3Xm1mtJeeeiKOuHldvXLxxMcdLuPs0TbGuEMc5cHmsIsyrEQCxJce9c3ciJgoRtsVnCABkSXTr3eoAWus4HJ4/fz4MQ6211qqt+exKjgb7zzagf25oGWrIDgzAAPdO4Z1HZ//Wb3z37/3tX/+NX/037l9cJGatlRgQ3E3dmrdaygRugBA1fAUfp7FpYyadPwVL7M7sPzE3a4x4cnLCSNZ8HMdxHEsppg3BmWW73XRdD44xLtK0mTZTTTlLSgjQdV3XdYgozCEAEhYCCP9zqaVOReNNCh5nJxQnpWltytFGd6/qFXhs7enV/lDMwcl1SjIlOmT7R/9oNXKsWbNmzZo1a76WFUCvWbNmzZo1a76WH/3O76A0QjBVIsiZz05OGA11ZCtW9t4GgsaEwswp19purq/qNJi2zAQAgJi7DgG0NZaESM3MHNS01sIEOXHfJURvtUgiInRHV1cFbWYG6uEmBox+LbEECSMBFJRMXQ+tojcEZ0JCt1YcwRmbtlLqNE2tqTkwC6WEkowSkABLFpYkJAnzpjrtrw+fP/nyo08e//BH77/3/sfvf/j5V88vn19eX17vgr0AooODOxMDRKt3GRR3qwV9W8WAMSHN7OLi4sGDB+++++6DBw8uLi6ij+wIh8Nhd7O7vroq02SqiGRmrVUANLegkGGimEcLWtMo57IEsQpMdqx/znRyqQnPpl+HaFPWWhEw9NzRo8VlfiAcZybCLOw47s78zHUWGSOTA6i2+MtjV5c5phdqcMx5qiHMxW1mnqYSSFG1Bd90N2va5S62Z+mfzlg8NszdkTk0F9H5jQJyYEp3j6ciomCPc88XEXEu6robsxDRsbkswoG2YzfjGUQ4DrKZqbYA0MEuVZWIRZjnLdF5FQCptfAUIywYNLwQweWTSLDG246OUKMsnWI0M1MPV3K8Yug1cs7BW6dSyjSlnJmJCI+slpnjmMeJCkBcayWJozGvgjDzy9/0j4Jvd4nzhPEMbsucyRnhIoR9W1+SaFdVAMw5L81uFJGcs6qrai0lALabRXH6ltcCYLkJAG4NTjy2dHGWxswQ/OjaPl7Yx8fHOyJq9XorcbhifKVZ3ByAzLIch1mTTfOkS1+uboibFlRnC0cZp3EchsP+MAzTNGorSAhIZrosWvx8GE3Lf1DRYgLZCJxt0v2752+8dvHuo1e+++1vvfX6w9deubvtsBNI2Miqt6kMe3Al9NbMkVCSmremrUzgjghIJDnlnK+vr6dxhFihEcm5E0mEYmbjOB0OB1qWBEQSINWm8R7vc2Yid5eciNHifaGq2tCNAIQlMQuzWnMwYamllGlkilMfsm9rZg6zP3tu0xM1kOJUjUf1BtgAjOTL03pnSp2m/+A//m/+337ErFmzZs2aNWv+BmYF0GvWrFmzZs2aOe7+1Wcf7C+vhhcH7qeOs5DnxB02KHvUguDWJq1FvQIYAaSua6Xsnn+lraBryimw4/b0NOYEIpGaT6U6kiNqa8wowjkJgjetUTmMG/WtmRkACXJWAEAiFhYRJgYQZuJkjk7sLFZG0IpobgrevBVzVddm2lprtaoDkOR+y7lH6Tx1lDvp+i4nRKrqX11Pnz158ZP3Pvjgg48+/OnHP/ngpx9/+uSzJ5fH0WPhlVgksz43KIOdzffpfw1KRXeViM7unJ+fnZ9st3fv3n3llVfefPPNi4uLnPPl5fXli8vnL55fXV3t93utDQCYKOfuaHJwt2maomQKS1l1qqVpc3MWDrVx1K+jFupHO0NYLxxmY4M5Ix/JIwAwzyMBjyiQFgezzhrfeV4Z3Op0x9dRzW5N49jES6vq4iae+S8zq1rIEyJhdl7sDg4AwXr7ricmbVFxn/8KfBFQuBEzLD4NADDT29eqqgZfhhmXL+be2TGipdTQV0fxGZFynu3SsSEh+ojyb5Dl1hqAxzhHAI+dJaKu69y9lBpFckQqtc62ZSKMI4aIiK01CF5P4O6lFAAgoqC30zS5WzTEVbXWqs2IFwCtqqrBEYm51lpLkZSI8CiduL2zuOBwM5umQswxFfB4lGLJYcaIqiFQTsw048UQPARopvn4IwCAqarOHepaSxyo0KrMl80MzT0cDQGg5yl5ALcryRBmmKW/f2sSI9ymzMHEW5uHOsYfeRaPxDBMjk79sdoczxO3FyynPqA2MctsuF4a/QgANp/x5bAAIUlQe8RaSrDXw+EwjmOto7mr6jiOdkvNcbwAj1/R/Pkw02cFEABCAIdtgnsn6Ze/+c47bzx648H9e+fp1bv9w3tnpx13pDodvBXX6g5AQjkzJzMfdwdEZ+HcdanLKaVYqUIkyYlTaDsEiQEw3muSO2JeetLQzBGQCfvcM7GacmIiUNMyTWUca5m0FmuNHAiRCMwMwVNKZhrzJ+OEgUPc/xHOG9NwdBASNoOpInYbTBtPaV+0AqupoaCxNW7D9jd/67f+/B88a9asWbNmzZq/AVkB9Jo1a9asWbMGAOAH3/tf7tx99Po3f+397/3TZn7adw/Oz1CncvPVzYvPt13q+066TR3HYb+73F3VOoF7l5MwoVufUxI212kcpjKmlDfbk5Ozs2iigqP0HacM4EAECPUwtFLUtJZiakxMDuRAxKnbpO0WJAFxkE9383GMgX9T0dpUzcp4MKvMBK7uSgTNWtUKBCmlTdfnrk9dz6nH1IH00G1AErIA0n4/fvnl89/53T/4nf/z93/v9/7g6bOr/aGaaVOrakcAvWAlmGmvf60vHBMIfwZA95vN+Z3z7373u9/97ne/80vfBoD9fv/ixYsnT5589tln11c3pdRAaTNaR0KAUoo7MHPOOWQLM1xbJs011apNl86v+SwKYOa4Wz/nTEwxYWwZx+dqijYLImqtbk5Eahr1WDePQX8hYAhvQzygtXas7ka3t9aKhHhsWDt0XbeoJKKmzrUWVe37XlWnaQqqXmtdjBkzKwzSak1FBBBMTW22Z8AsNRZ3L1NBJiAEgKDkAEf8Ovd847DfYtAYld4oj0/TFNsWdNXnUXiSUgqqmHMuZYq+edf1seVx8HPORBTHAQA2m01rbb/fh0ol5253s5tKOTs76/teRK4uL809hhlG5dxM3VV1Rv993yEeVSGYc3KH1tpwGMw8Wta4eJ/dHWe5NrlZnO4ZTFOU5VutJU4QEZl5KSUoYex7NMejp+zxtMu+dCmFdtnd1MxUaS6SQy1VtRFzKDW22xN3Pxz2SyuZY7Wilrq079kdYhZonOJaSm2t7/so3iLR3ApHZJ4nIoZ+JKWUc46rbqljA8yg3eKacYejiTr2Omq5x4I1IpZSWmvzeyrK4cRE3GprrYXWJnq+ADD3o4WTSMxmJKYwQQNATmm76d29aau1HA6H3c3Ni8sX0Wr/el6+9Y8AOv5sgMsHhwtAItwwb4Q2id58ePLdb7/xb/+bv/r2o1dfvXOSodXhZtzfSLyzmPt+wyTlMDgAC/fbbZxujOGKzJISCTtCrVqKAmC/2ZydnWPOten+6kpVESl1HZNwuDJqG4eBJBZrsNVapnEaxmkcpnHwpqqttsJIMVw0rplbfpv4DCZzczM37XPebvpaq5o7sDo2kEZJtmfK9GI3FlX1Mn71SuqvRPZ//x+vOo41a9asWbNmzQqg16xZs2bNmr/x+d73vpfhINjAi1DqM283mw48TXtpg037abjCkBsQl1LHaSpaAUESSxZmjjl14FBbczNA7Lsu933ue9PmAMBC4GBaS52LizV0q+4AhCgkHE8ETgCIYOCttmkqUZP0ub6JBmKAFgCIkYQBARlz7oDQY5KdiOSOiRHQ1Sj1lHpHfn518/iLL3/wo/c++uSzL7+6eu/9Tz748NPPv3g6jKWpH8fazf+b+dL8yxLi0aR7S/e8mDfu3r376NGjt95669VXXz09P4sGK7jvbnZX11fjME7TOE2lVUXAlNLMZN0IiRDV1B0QgFlwaTEfzRLu7ggzUF5G5yHBseo6Ezr3UgsgBquKe+dBgYkl/T/svduvJceV5rcuEZG597nUhcU7WWSJpKjpprrdbrchewDb8zoYowE/6J+wYdiGHzyYl/4HbMMw7AGMefaDjMFgYHiM8U3j8aDV7unWtCyJakm8SaREssiqOnUue2dGxFrLDysizymSsoSewbhJ5QdKVWefvTNzZ0buc+qLL35fKKV4X5xvb4lIAwIhIXm3oTpB29SqVM+QOg6ilOJdhIuZ66lnEUkpImKt4v7mdrvxzr0YPT9bFmrzksUmREYSETV1NohzKapUEYkhIiECOpUDCbGjGJybvHCWHX8s4vQPEmlY5CXBvfAuloSsFx92RkdDK7gH6rCXxd18NDnuwXBrprBhzllVh2EgIvAzDxBjS/66ke20ioZ76P6479d9diKa5+JvJ8XoKXhHbTS4NpF3FnpBn4MylvpEv/odD1LVFBA5BO0FiW4mVhHpUxpmxl7H55WZbfw40qQAIgJ685yZOSx4QX84i9rAHNgzE7/9AAAgAElEQVTNTN4lmHP2tKyZ+Y6I2U9Ce6cxLgPZISrLCWl3d0/GQ7vv7Gpi2u8zDz33a0qLB+0rKLjhR1BVfabKvX+/+oTExJ55J26Rd1UFU58V8KFLxDGwmvb8L5jqPM/zNE3zPE37Wmp/I+rNo3jpPEMvJ7xcKEFgBBAAAkJAODyIj904evbpx1946vqdZx57+fYzzz/92NOPX0sMaFVqDkwIWLNQIA7BQ+VS6xBi4EBEaqYqopJzKblNMAxpFDAHuJiqgTGyqqk4NNzPORIhE4uId0KK6lKeWWvtIXUMHJi5Sq9kbHa610siqCACkw9pQmJRqApFAcdDjONc5MHDhyfn5/tdQdjXWqtUK/uv/8H/8Bf/EbVq1apVq1at+vxrNaBXrVq1atWqX2v9+I/+QcFhx9eO4F4IISXebNM2sZ3ekwcfsQppRSu9EQ2KgiBgiCGFmAJFRGZgFgMRzVkCO7Y0MZMhWi0GBjFAzjJN8zTVUkWt5W4RPbgYyLEAIKVYzVCzlDxP0+7iPIQYQkAOaqRAxAk4QgicIqWIMQARBh7SSCEAkwEaMXBAA611vtgXgSy6O9u/9ZP3vvv6j/+vb/3fP3rrJw/P9qdn035fLvGu/dciw25AX4k3Yw9Dm7qbQyGEzWaz3W4PDg6eeeaZO3fuvPDCCzcfuxlTunv37vsffPDhhx+enJxcXFw4gWEcx0iRiTsR2HLJ3epCU2v+GiCYheCZ4nbmkamVKy4VggRuonn2042eXCoHZmbqph4CMnIIwTeFl6Y14FUfEwEBDcxNagAwcFRsyymLiPfEeeWgO55ubKWUEGGaWl/cMAxuszIzgJXi6VR227eUCgCBOYXoHi61ALVPYBQHNAcOMcU5F0+wAoCqlFJijMMw5py9XG4YBkTKefYrUqv3DZIHWsdxdC7wJYOhG8oO3Z5nrzcMOedai6qmNPj0QCml523BX9jz6WRm81x8j8wstZZSrhjXAABm0C5cf8h6HaUfg4h4BFgVWob9igEt3YD2FLYb0Mt5cA99ccmZyXfXSBdE2ujV5KHp1rDX3VvQBt0m9Jh122zOJaXIHOZ5aulgaqa8W8kO1tBmXHpgfwTAeZp8v2Cm3bX30kZRZaJxuzWwWqsPhpQuEdvDMPjoNXN6R7eizfz4l8y4tnpA6G+/nVVEQiCidoNIbWxoa8WG2EY3kJmpdZAOtOkq6Lv0eRefdUCEGOMwDkNKCFBy3u/3FxcXOecqUkqpUlSbabtA4dsNdYnj8AcNAQiArnzryZvbO8/e/Fd+49Xf+eorv/0bX7pxmMZgKBOZgqmKxSHGGEqtpRStMoYYyE++1FpLKTnnWso4jERkaqUWNE0x+joBU6211FIRwe8vUEBAIhIzM+AQKQQgRkI1ENHF8SdiACylmBl1ULiTyon8I8JHIxExI4qBqFWxaijInLZTnu+fnDw4PS1VZ1Xd3Q/j9RiO/93/9D//C/+cWrVq1apVq1Z93rUa0KtWrVq1atWvqT74zj8UQTGbiwBiHOLNm1vTOl/cz7tT2F/gfifzjKox4DgMISakwOOGxi2OAyCQCpACIQQGDobBFEENVVGk5jzPc81ZpQKp1Cq1mhozxRBTSDHGEGJbYw8gpeR5Pj87RZPEaLXWMpd5HsfNMG7iuMUQjdiqYEi42WKKECPEANDork6FLaVWATUMaSNqDx+e/fS9n7399k9//KM3//xHP/3hmz+7f35+MeeqDU0Mnlv8Rb8TmcN2AQkI3elTANhsNrdu3Xr11Ve//OUvP/fcc5vNRkTefffd+w/u76fpYrfLOSMAdsqtW2GMwdQc8ezZ0mZTEopInnOLZyIOaQghTNPUssZmC0jXTWrrmJDuvbYALBER83L4iRMCqmktjbDhj6tpTw3LJ5LOV/O5/lp/pNTqxqj3zDnWmQjdDO35Vn+Q3Kh1W6+bv360gEgE6Ba51x66UZtSAgNRcRM8hLCbpirVrVgz2+/3zJTS4IWN8zxvt9sY434/OeV5GEZEcIeOiDab7TRNtdZhGIhQ1RwSYgYxBjObpimlwXHMIlVEgndiIs7zLFKJnKAtiOhthP5Gcq4xxhgjE1WRUrKZm64teb2Eqd1kd/fWE9Aex3Z3m5gCR68Q7CgUEhEVUTNPjrdIL9oSIfcJgFIqEfpmzUzEJ0bwEwJoJySXMg7DOI5M3gZZPSnvqW3/R4Gb7/7eVc1d72EY/NqllGotnUfhG0dT80N1K3ZpGPSIbMM4IMIV1vPCjSmlbDabPjvi3vUjhOiejwYR8c8JjyovmBERQaAO7wYkjDGa2jRNDhIRVUJEQneJsZdnMjNdWefgrndjWHfQNvTzEkOI0dss6zTPp6cPz87Pp2mPrY2zLGn05SXLTMRl72H/fwIMAYcUjjfj7aeuvfLCY7/56osvPnPrievbxECgVvOQYkpJRVTEVK0qmBFijJGYaynznEuuB9utmc3TXqQCGBMOMQXm1lAKGFNypvzyAWcKqqCAwEQh5FprFRUNQ/TrgkBgWGtBpBSjqgACc1imZJiIAoqIipppqzs1VEAFUGQ1rqI8jkVsVlOyZFsMFVER4a//h//1r/TzadWqVatWrVr1xdJqQK9atWrVqlW/jnrrj/43DjpEK4UwWWQMhKDTvDvJ01ktU0IcmE2UOcRxTGngEBGQQ6IYIQQwA60g2bQKiBmagilIrVIqmGqVIlVFDBSos3sJGYmRhhiZmZCqaq3SqMO1llyIMAXHoiIyhTTENHBMSARgJhXAkKhUpx2zGpgvuydColxsLjBnuH+2e/+j+2+89dM33/7JW++8+/P37969++DjB2cVQB2osVAI8DLrvACelwdauBEhxXR4eOS9go899tjNmzdv3LhxdHTEzLvd7uTk5N69e2fnZ7mU3W5XRYaUsNnryEwhBBWoteacYwhEPOcZrVWxqWou2T1I6HnDZlMSZfeFydPShIhq4gxoWMDBABz4CqQaEaCVEEpbTc/EanqVUHH17wCw7NGPBK94mkVEVT3L7C90p/WSE9IDqtBdN4cdiIg7mH5aQwgNjdLdeYcetCg0Ui8JtKqij1h7tmzWKR8pJbdo3bWMMXlzoLv2zKGUXKtnh82TqosbqKqlVKdxe/RbpIYYCElNaymi6ha8c6U90EpIAFirNI4KQL2kbTziQjIHZu6HpguBYpl7cGs+pcH9aD91IQQE8Po7vxDYugTJrJ3phknu2BA/A/OckRCZQ0dpM7P15kZVq7UOKQ0pEZKqXi1gdE+W6JL37ShsAwscxnF0495p7B4G90hyreLzDSEEwka96IMPfRLCFihFd3UXJ90bF5tzbZf8jcXPXdLrquZDcqFz+BZqrURMyJ3lQiEE8Hh+CzUvZx4Q27lCxBijSFVPhXfOtKlKFe4DX0RVxUwDs1/uluPOZZrn3e5iv99N+33OsyxX36k8fbhCf+jqZ8vyr69AcLyNN4/H5596/Olbx0/cGG4/9dhTN4+OBx4DJfbryT5hAAZEaAZqWqsAIFGIKanqPE0xRmJCM2YObT2BLa66TzYAQHeNgUMEJAWd51lEmBAJwJstAdGwDw9uXBSwUqtUQaQQAkeupdRO81jelhqoIQASh+HwGnIqJmKohGBKaGd1OJP03kX6g7WccNWqVatWrfo102pAr1q1atWqVb9eevub37RBjAwBMdoQ7fhwGzRP53fvffiuaAUEZD48ODg6OiIOYdjG7REgGwCIgniCzsDUTGzaybwreZJStFQT9aAcBUJmCIEIgQmYY4ohBiZWERMdQkAwFZln7wAr5nyHOHCIgTgNQxzHuN0CsQOYTYpJNitQM+V5f3ZWcgHmqqDAIQ0hDRTjftKzvTw4r6//+J3vvP7GP/2z77/z7s/v3jup2pbAd/e5IVvxym9D2PxmgPYEQEQM7J1pR0dHzzzzzEsvvfTyyy8/9dRTKaWTk5O7d+++++67H3744f379zebTYgRCX21fhoGN9aZOQ3DOAylSCm1Sk0xMXPOORA7e8GtusbB8No5M4drE9Kc5+ZItjo+8AR0jNHMci4AhoQUgvUQag+oNuCCO2jEjnRoLI6FC+GsgwZo9vxyCyxjiME9U09Khw7bNVMkiiHU6riF6q8dx0FEc869F4483xpCcC92GBICSBUmBgTfkZmJSgghxVSleoMchQAIywFvtxuvN4wxdiaDIWKMwQAcWeuWY89ct5S7iIpWM02dvu0QDwByd80RKKoaIqPzRroJ6hwMH9UiEoNTOICZELFWPyvqEANHRXsemYi8Fc8DvO70AZiHrLtnDTEOiGSqVQQRh5S80M/PJwAwEQcKgbVbim7q+gEAgJ/YaZoAkUJIMbrhGlMys1pLCJGw0VqICPTSI4ZmxGft2XYHJbcWSsLAIaU0Tft5nmsVn0cJITqDpZRqaks7Yq0Vuju8GNCA2IDjdjXE3eTuvDvARNTnPtqB5ZzhkuVNRBRjM6yXWQdCdlAI9lvDLXuP/ONl8SP5gPQ5gBhjztmT8sxtC6YqpaYYudviDj/pcw/t/huGgRD3+/39+/fu3783TbviV7MhPJaPk/635RPmUaQPM4IBqAWAbYLjLfzub7782kvPvnjr6DjhyLjdbjfjOAxDW9zANE/TPM8iNmw24/bQAKpoKfXo6DCmJH0aI4akqjmXnGcTJULmAAi+5AIMttstmJWcp2mPoJsx5TKL1MCMQIvZbWrEZGC5lBbER+TAxI0lXcQT0Asf3wwgcIwxCaAhG/FweE3A9lM2KRjDtz48vHN0djRM/95/8N/8RX+IrVq1atWqVas+f1oN6FWrVq1aterXSG985x/yTHAR9FoBs6ODGNHk4gGUHeqEVnhIPA4QYhiGMAxQDQ2JohbRUmupYIYGpiZSpZSL85M8XUjJoEJmEYkZQ+TNZhM2A4wDtrI8BDTPddZcpEoKEQFNxEwNDIA4DZxGHDcIhKrEwa0sEc1VpnnO0/m8P592p5HsYDOAGnMaNwdzFkE+uvVEzuX+vQev/+itP3/j3R+++bO3f3b/vbsnHz88u5jmnAsRGYCaGlLnbvxyAzqEcHjt+Pnnn79z587t27evXbvmZIzT09OPP/54nme36ryozHHJRQQBiZCYa61SZRgSIqoZAnlxX+gyVa3ij4zj6N6fs4lTSqICS764RSxbCLYHQkFFqkgIjESAKK3ksUdHa/WMszf7qapUMbMQg6p6QyAigkEpRU1TSstz3P5uNFgisWZPQ6cfACBxO4Z5ziFwjMm97Jxn9ivYQ9bu/bltTYBozXR2GrKDmxGRiZHQzKQKeOVdD2Wn5L6nx2ahx4rBt4mIKgIADmRAxGEYSim1luWKeihWREqtYBZiRMeqVIkxpBRLbUbzMAxMtNTreSq5u7TsMVyncxARczDTK+4i+Dlx5kmzOMnB383nXai7PStMJWcAiCldTaNLrT6ozFRNsVUOOsuikR48HC0i2HfmB8DMalpKQUA1c3fSzFTEp2KiG+TM85xVlbklo5dA/OJ411prFbdunUPi9nzJpTnvPQHtp8u95u4p+w2tCxu6VnEfuQeUfVw5utwxJLRYzL6FUgoRxxj8wVKKR7xjjI7N8DFs5kQQLwdEvPKHX+iFyr0E4S9NfTP/nHLwxyU/BC7J6764gIOnjFlVqpRS8n6/3+0ucs4lzznn5WbtrYRXPl6WWS8/LAMAY4BAFhFuHh48eW188Ub4yotPf+WlF15+6UuHB1swQRNmTDHGQF68SRwxxFykiojCMA5+qzIRMyMSmKlodcw6oZkagn9EICAhoCmaqgiiBWYf4KYNhN2Gkk8RGZh5uhnAUE2qCnEgDj7yVVQ6vcSBJ4AoamqARBAHIyqip+dnFxfzrkx7qyFkDXM+3n/962s54apVq1atWvVrofD/9wGsWrVq1apVq/5lyL7xjfvX43Se94cppZIixpi2AXA+y7rDIMwxxQ2nyCE6SQFFNBfJUqpqrlLEA3QiWrziLAYBw5hCYEJgxMgUYogpDOMQIkMLlppWFVVRqaKOHFVGpkAxEBMSEhKHSCEqB6lV8lwxu0M57ec5l2pqVsEghEgEyjFtxjQcpO3xw48fPDg5/2B394P37775xtvf/9E7b7zzs3fe/fDe6Xy2Lw7cQCRAArArsGf7xJ9t6TyCmaU0HB8d33r81q3Hbl27fv2JJ5988sknDw4OVOT84vzk5OTBgwf37t0HAGIi4hDTlkMMQc0ozyFGJjZTS2YtTugFaAwAIuLGX4xBRSsVrMjMHAJIJaMQI4fgeIVmw3WQdFUBVSJyZHCtFdCDrYSICoBoRJdte9rMMDQ0M8ilgBki+bdE1d1VN5Hcb1O1qgIAZARm3omXYrTWPeiL7r0yrtE8zBqY2Fm0/mCtxW3KJUTcoNUe/RXzrHcD/iJ5013F6maimi41kG5WTlOLlEpb+G/9f80vU/FMtCIYAqpUBGOmq4WLvtlghojDOFL3JZk5psCZhIOBDWloBpwTMIj9aJ3zwBQ8yeuWtKM/PG7tR8stNF0AvK+SQ4h+5H6lCFtit7qBS2QhXPFC2zD1Nw4GZuoeqEJjSkj10QriAAlCUz8BHvT3FkSRKn5gLdZt3SpH0D4Oc84iyj0d74OLiQywDQxruWuRtvd2ITpapdbaGiwJmbjNDQA4sMXvKfea/QOks7CbVJVJTb1ZsRmgHrJ2x79hTFRE7TL7TOTVgr7Btm6g389+komJiYnIQFUaqcZUVc2HpR9nQz9bI1tfjei09RJwydLAgkzE7kP7511MMcZa6zxPF7tdmXMpxXo5IVgbfs7BsJaMNp/LQwNBMIFq8MH9i9PTiwf34GSyjyf+aKann7h542h7bZOOxohABBgJh2EAYlE0tBADx1RFpGaTCsAIPv6BzQIpkBFa1qpmiBRCDEwiBVTIBMgteuMQEbHNCPm0CrFTXDzWbdAmS0SlSqEQOcQYon/CVxETn6JAQFAwEaci0ZR31eDg4HhI1zfp9P6J0gy6l7Nn9/jxtW/8F//x1/+T//JX+RG2atWqVatWrfpca01Ar1q1atWqVV98/fk/+fvXZnnqXn3zzpYCXTveHgwx2b7sTtEkMsEYITAYQClWSt3vQQ3NyjSVKZdpNgUVq1J303wxz7s8b4+Pbz3x5MHxQdqMoUUpCcggEDABGkwTXFxIKXXOeVeqqAJYIAU0wO14MAybNAyQAiCCZBAz0TLP0+5iv9upVgAkiienZ3Mp2+PDw+Pjw+PDYRzUdMp5e3gcxyOIB3/++o9e/94P33zr3X/2Z9//9ne+/9Fp3s0CAAqgnmNGgoVIa/aJSPEiz/Z6YvfGjRuvvPLK1772tddee+1gezTP84MHD958880PPvjg5OGJr+VPKYUYANEDpIg4jiMATNPksNpSioOA9/s9Ii7NaR6bdSfW7UKR6svbHbzgbWAAMKRRVD1T6TZlLsVUh2Fw/27O2Y/ceh6YCMx0nrO7hAtcmJnNdJpmP3giFE9AE2PzB9UMHHS7tMAx8X6/B4DNZuN8CQ+fErFzErw7DhEdBOGkYKdDTNPkX242GyLa7XaI4HtX0TzNtPjmbhwTdu6B+PlUM+qtg94T6BjfUorv1BPTMQQHlXgAVlU3mxERpmnyqsDmcoI53QJ8DoBoHEfPIBORmooIGjCRXylPo185e6aqHtMeh22ttUoFgBBCDBERPZkLHWmSSy65XB1gyxMWmUFp/OWeK+8gEXMIrzOLwZiaE+1GbAettBHMzDHFKlUNPNLuw8xjxy0S30gXtKC3e9IX5zmLiBvQquoGNEILU6vIgqRQVVP1W0lUkekqzsJ6x6BTWUSqQ7rdIAcAkQpXgONXDGgLPqQQfUmBX5ppmlJKTjr2ZD9xcArNfr9Xs34F3ZX2+QBuuXtRAGhw5J7Edw+6oWY4EDF1LDV0ljqAM98/kWi/8kEBCF4jyRRi3Gw2ITAREFHO+ezs7OHJw4vzcynZywABvPlTQ2BA8OUFAACEbRBYC0cTAPV/nqVIz9yMr71y+/d++ze+/NStZ24cXt9EKReMcuPmdUSqRXKVMIyHx9fvP3iw2+/QNBAGRCIjUzKLgZkQAGapXng6juMwpCpFa9Y6mxEgI8aYNiEkv8FL9Y+FJlHNc0Ek5uCLD8xUwQCJicHQp3BUFZoBjeYTTAhMtNvvi8rm8DCkEYnnkt//6MH987kqVN4EE2b8/f/ov/olP8NWrVq1atWqVZ9zrQb0qlWrVq1a9UWWfeMbD67zPtFZoCHaZjscHh/GCEH2VHdaC4igmhKIWS1SSqm5SCklz5IzApIaqYICE6VhhJQ0BCEIm81weBACMSKa+vJsMym1ZM9+1gKlmqhVA7E0DHEYMEVghhCYEgORyD5PU5lLnn1dutRay1zzjGDDOF47vlZUKxjHGDfbOG6Qg6jNVdTo3oOzH77xk2/94be/850fnjy8uHvv5O69k6loVYC2+h0uo6Q9cQmestTLBj/opW2PP/74Cy+8cOfOnaeffvr69euIKFX2++n07Ozs9Gye53mec85VqhvKxGwAbkqGENwpZidviHSTdCl5a3+JMbrV5YhbT2I68daNSGiEDSZsNrH71J6kdvPK49odtUFeU8YO3YaWU3acsb82xuiFgeghXmp2LTd4LvRfCzucAMHtzuZ9N+vWahX/Erph18EP5KCGToTQRghRTSk5YQP6pfBdLhuH5ssrEQUOoiJVSi1IFGIchkFEai1OWsCGGIY2o6DmSd7AARHVVEXdRi+lxBiYWUWrSisVJCTEBhpY4saIIlJLNVUEZG6ID5G6mLxL5BkAmKIHRQHAg6LubaqoNz2GEC7dzK7FeL0qscbggE8b0NQuEyHGQJcwFmclqAF6KSL4coRSq4GF4ETshlqm1rAHHTgB1gDN2C1fzDmbwTAkaYWKhtjS3767YRh8VKuqAQRm8MuHrVvU494dOcJLVWC3whuKZBmuqtLbARtHBQG8cw+Xs+20kH7i2syEARIHZq/lTCktPnY74eadjdxw6qLW7Glh5iENzvsutZj1FlJ7RD7OHZ3RLw0uT+qfLO2ThJicLaMiwzAgYSnF1Gqt8363u9jt95O2jlRFNCeF+L3myfZlGgz7bY1ggMiEBwPeOjp4+sa1Z47H27cOv/TszeefvfX4zeMQoM0AiCARx+H8/KzWklJkAkYAUFRFUyYk3yNSVZvLHGIchoQICIomoiaKKgwUANsVF9H9fm9mPrGIgKqGyG3lhNYqWVWRKHByz9wHlkONAG0xoKm1xarfyyENnMYseDZVRVILFHmogUsM8/jX1mbCVatWrVq16our1YBetWrVqlWrvrB6+5t/b8z61EN5+86ACjHhjaPDzYBYHlqdrMxS1URBzRkb85xL1aqGCFKrSB1iihwCEQAEDtvNJo4jDdEQgMkCgorVqrVqraaqYPM0T1NrzAscwACNGGl7cDBsN0RohAYoYlYqlny2uzjbXVzs9yGkNAwcApqCCgXabMfrx0dAqIgKQGnEOO5nPTnb3Xtweu/+6Vtvv/cn3/7en3779TfeeLcoFAVpacLLcPOC3Gg0gytpx2UN/rVr127evHl8fPzUU0/dvn3bWc9m9v7777///vv3H5ycnp7td/txHJkZwEqpZsrMSOQGNDOnlC4uLlQlhNiTpC1z7dlhVfNEbUxRRWunMy8BW5FKxG59OhvB7WM31zxOCIBeagdg4DYikmeowfOehNAMI/Cd+jM9o45EThNw/sMi6CFcVVnyqot1eHVQtS5Eah5iP40Lz9cQwbOo7juLSD8k7a2HwESBO6jBzN3teZ4JiQMTNjseCDkEx1IvTzazJcmr6hMWhRA96LpkhEWa5+hXIZdSarnydkFUSi5qbfrBab4qAoCL96rqBrQ1BES3y8HQ9+LnzQ/4qinsBj10u9n/ICIOAa7+/o3d46TLE37lm+Qxc2ZKIbS2N+sY8Mb64HYMTFXEDWhwoK8oEbXyyeZlL2yMNg+xRIMRcRiGWqtjdoiYObSRZzakxCFoB3D4Lpp53EP9Plb9zfgMig9g36UfwzJ4ahWP/1/avtCOxgeqg1+ggUR08bJFW1mpiCJCZ0DLct60TSEwMTWyuaqolFJCCJtx4/dazrnjSrorD91WXqxh6F42oqPG2/BdcN/obI0WlvdmUUCIMRJSnufdbre72Jcyl1qkZpGW3PdXmdqC9bgyKNAZ0YRIoNEgARxHeOrG5uXnbr368nO3n721HcLxZjgaEzd6jpSaASwNyePgZoZghEBtsk2R2AyKVGIOkZmQyN1wVMVaURRU/XMAAXC3uxDVQAxtvsrdZwIwkVzKpCqAFDg1dDYAARKCmvi7Up8zYyfvO6McmAPGGMZDCgPGzVxVVaDQcHpNDk55O/21f/+//cyfZatWrVq1atWqz7tWA3rVqlWrVq36AsrMPvrJ6/nhx+X+/RxxTHZ8MBwGxHyG+Qw1S8k152nKYogcZ9G56jwXoMBp2Gy3w2ZM4ziMiVPCNLhri6pYi+W9Xpxbnc2qqkotc87SLNJYxKoYhTRutgeHR0hMSITAm5FigP1e9vuy2+0vzlQqMV3M5Wy/f3B+cXB87drNx67fuD4MiQloiERAVkrJtRY1COMBhM0Hd89e/9Hbf/LPvvf66z96482fv/fzh7v9PJdavSMMQdyJ+lTUFNrDLW3qXrBX//3O7/zO1772tVdffTWEcO/evZ///Of37t3bNe13+2nOudbCHNzIwyUV26DJ2sgSqrXWaZr8S086q2pK0ffoPqaomBoRbbdb6BZbCGG7Hd3m7MhZK7l4s59naUOIXkbX85cQQsBWv9a61/rbJGvbabVuph3fawCG1mkJzr/1IDMAOObCw6qLh3hpvPbAuJmVkh3ZQYSqOk1TSkNKyfPa3VYlpz+riruWzd02M1U/eBUdx5GYLi4uPD263W6bS1iLqCBiSimE2LAOtXZqAnrSXOLyAbQAACAASURBVEqRKlXqst+5lJJLLtX5Gh5On6ZpAZX4G5EqntXlwKpai3gW12PFAKZawTnL4rjj5pU7RnlxgRERu31vHSXsp30ZdZ/4y0J+wNCA3nCJZ2FqVXIIgMzERN0KxKsb8dz3MqrFFBCYw7IpJ5aEELzfzwcJEWojeKhPGwzDEAKbQc6trtMNaPemaynuQbbOTFWvGRQR6BMPjWvdbeJaG47DvWOfTQGAUko/AM9SXxrQgZmJa61ElGIUVW3hfTAAb6qMMSmAapvrYOY0JFUtpeZ5DiEM4+C3pbvkiCjN5oY+jMFRLbVWXI65jUo001rFTXc3tdEXOhAhkp8x377ntQ0bkNsh47VUEVEz7xd1zx0Azs9Pz87Ozs5Op91FzfnK7Njlx9IjXxEiGAGwKQGQASEkwoPIN4/jM08cv/bKnddeeeErLz5zNEayUqazGAMRK2IRqSKAyCHEmIgI1KpUrYpAwzggOkZcAA0ZYxyIWBRqUYeWBOYYAjH7WZrn2dRCSN4tGCKbVZFZRMwA0XErhkAxcAy8GNCtgpAa9EZNRatoBSLAoMgUNwJ0vtvtd/syy2aUaS95lt//W3/nMz+6V61atWrVqlWfa60G9KpVq1atWvVF0/e+941r43PPvfRv/OAf/90x4WYTN4GDFZoeyO5M5gutGdxSRCJOFIdiKEjAEYaR0xhjDDFyZDZT02rga8xlnlkrabV5L3mqeTarIrVWoRBCGtLmwDgaBRw2IQ6JgxmaaZXs8VfMxfIs817yBKAcglGoQJNZOjgcj47GcQhMCDDXolq5ZYhBAD++f/rOex/+8Z/84PUf/fSdn3zw/of37j84u7iobgtZs7+gil01TD8tNzQPDg6+9KUv3b59++bNm0888cTNmzdV9ezs7O7duycnJ+fn5zlnJ9tWNYceIzRTVUXMw8vMBlBrRUQ3vMy0lOqAiLY2Xz0x2iDLbkB7SNPxxB3QgSEEa8xqgsaWECYKMaq0uLFze7VnWXsmWntOEx394d6fO+PuCZZS1JSITGHZlD/NfcmuVrfmUOAYo8e9F4CD+7NuK5tpX5UvIhJCYA7eR+cerqMetNOl3XAMIYI1bgZfMVu9/8zUiClwYOa55FKLqjIHZhLRUkrOubEgevBWRbWKaMMvENGcS6ni+AU3QKVKLtk9TYNmMTe3H5CZVEWk+O/GuBASvC+um6TQc+KftBC7Nezus4Et8eLLZ1w5vXDVkm5lhNR31CAVxOyvCoEZaTFJr8qH0HIIQIiEVwzoZv72PYI1Z9xXAPR4c4snt0EiojFG5kDUCjPdFHZ0tE+QMDP49pnUoJTSEPDQONG+C+jTFdQj3iJyhSTziAgJAWqthH4jQDvbyxNahD8YgIpYx+a0okUzT8E3rPMyEwPoFYgehTYDZiIk6MWUl9cC0SEr0OoGL9Er/dS3bXK3rTvep90RIlJFfKaKmRHBD6ZKqbXUWss8z/M87Xf7/ZTz7NV+j/5z7HL9BgEQ2EKiJgQ2GCNc26Znbz328nM3X7l96+Xnn37+qceeunUcmRCsiPj49/5SpIALytyQkVNKbgQDqO+gXWU1E1MxAGDvnzQjpBDCPM+iQhS8bNBMRbNpJmbiwBScL9K5QLacV1UFRKagl2gOAIRSqwEiBQqR0saITh8+fHDy4PxiqrOQRNJxC9dWHMeqVatWrVr1BdNqQK9atWrVqlVfKP3wm/+9JNRrzPeAgx1sN7eONrY/K6d35/MHMs9SZlHhGFMah80mpjHEoRpijHG7hWFjIZkHOVVtnmue53k2VSm1zHNkDExoUksu8wxQDRQA0jAOm4PNwSGnEUKyNJqBlapVSi1zmUopWoUU0ARNGIUJmTltDsIwYkqQkgV2b1cV9tMsqhx4znU/l/P9/IMfvvVP//S7//s/+uOf/PSj3QRVQQ2wg56JyFfEV1FHyn5CHoochmGz2Vy/fv2JJ5783d/9V7/yla/cuHFjv99//PHHb7751kcf3T07O/MV97q04RGlYUgpecSYiEou6uxjZgO4gnJuzqDnKN2A9iio28QeTF7oH9pkTmcWqUtweCEcuBvpacSc58CBOmRZVRHMDNQsxUjEZuDmLCJ6hNOBvKriweQQghk4nmLBLwAYElm358zpsrUZ0J47bs5qRx4vCA4PUC9MDwBQU4QGaIYezvXvutkdQnRygJtcMUaPhDd2hGopBQlTSpNPANTqF3AxoK940Gp6GQrvYWQsReTSSWz0FTVpbYcIRAEXoLYBIplW1QJ41V+2SyN6QWNf0aXpfGlIf8YTPjEIPzUwFRD7fg08Y4uISI4K5hAI0NS6+3yZNvak7bJlYnc+vSbOut3chtnC/nan+IrBCj0X7qlkGIbEHBDaC0U1hEBE0n1/Zna7lkMwg1KKVxuCQZXq9BXPti/YakdRLwiOxeG9BJsYgIMa3KIG8M675Z34OOMQG366b0FETZW6J87eSEk+E2NMjEQANs+zSHPDQ+B2b+pypZdrcyXVjgh9qYRPPvkjTK3x0nHmxA7CIXd7c8lLYhoACDFEXw8RzCzP+ez09Ozs7OLiopZZRR8ZEWie3/aBR/2AsOPZCSAAjACPHYVnH9/89qsv/dZfeem3/8qXDjdpCARShyGMKXrgHbDhenKpgULgGAKLSJUKZECGBO0Cqzb32Eew2jTPIYSD7UGVKqIGIFVqqblkkQJQ0jDEmJgCESOQGkitohVb42K7bYi4X2LwUbSfZgOIcQBE5BCGVEUfnpx8+NGD3VRyxcfg9p7vayh/42/+7U/dLKtWrVq1atWqz6tWA3rVqlWrVq36guib3/zmsZ0nyAlnNUgRr984GMFgelguTvL+LO8uEDHENB4eps0BjxsaBiRCNZMKqgAmalWkzLnmIrkQqDditfQaYEgppKSAhkiEIRIFAiYkJmbyralJrSWXkrO2hesKSIAEwBwoBkqJvG+MUkJkqEVrqSXvpqmIKYXDJ5+juJ3O83e+94M/++7r3/n+62++9eF7P3tw/+R0motqA7EigjXzqv1W051CAujM1nbweuvW4y++eOerX/3qiy++8Nhjj+330/n5+enp6cOTk4enp3nO3adDA6u1ErGbv9QIG9IDntTNKRERz5Zagx5gjHGaJhFNKYnUUmqMTjMw56suAe1SWrFeCGFJj3bKASKCdUKxGbozuxh2fgxuKxNiiAEAvSEQAFTF/U+pYqbQDHrQBijpnqyHVS+NVGhWIAB1Nx16iLKnYNsLPdbdSwjZoRkd/huc3QFgROwY4h64VTPwgjk3l90o9HfnceZedmduQC/2KMBynrV/eaXG7YpFvHA2oD/WyL79wavZZGe3GGgzf6+Ys/DIpj+hT4aaP+sJv8Jv2rjs9BObuprPRa/Euwz2LgSPKx43tuvAIbDjYnybfoFCYP+2g8KXiYEOxGgupCfxwaCHxQF6ur/kXGsV1b5+ou3wcirF2qzJ0peI6KBk6jH83Ae/T7RgrdXMhmHwoPLi6fsKA0B0HIQHsUUEkbUtJujecb/YHogmN4I7r9khJIjgQX532xExxVhFrrZEop9V9AHmLJTLAQ8GxOS76wPSkBZDHxwtAlfi8o466RMeFAIvxA8RmfN8dno67fdlnheWdIf6XJmKWCLz/T8nMQ8BN5GON5unHtvefurod37zyy8/99SNkY8GGhmszpEpxmgIpUrOmSmFkEIMgGCq1SoxxEhznlQUgUOITAGwG815BoAQYwzRZw5KEZ9XQ1QkY/a5kNDnmFhFa5Vpzkvnql9MH3gOplexXCoAc0h+txsqxYgUGeF8yhezGnGI40MN55ber0d/sEahV61atWrVqi+EVgN61apVq1at+iLo53/yPz6Y4W4+fE4/NDQOdRjiQbRQLyjvJE9Si1allMK4GQ6POCbiIIgqorWYVFABs1pKKWXe76EqAaTQMAnNPibiOFAajAOESDF6FFLMucYK/p+IlKIiquIupnN2MQSgSIFDZGQzE5UqqlKqzjPUCmrAoRrNxjoe371//vr33/r2d3743T9/4613fnL/we5iV3SxaMBdp7aK/TKH6t4akFqDF1+/fv3xx5947rlnn3vu+WeffXYYBkTMOd+/f//hw4e7i91+2uecm+UK2MrlkJq16SYWc63FWcDuI7v9qmopRTOrVTwsyUy1VjMIIVxlFkN3daEZiFZKVTVE8qSnI6LhihfWzS8DXCzvqh4jZSbE4nt0ynPvDESAelkV6HnkRpUQ0W6rgVuGITAiXuYwO2TDAda1Voc8lFIWP86z4TEGjzm3WG6neTSiBJF1P9cPrAOcHZohWiUXZ5wUz0P76W1BZVVVrX5+W9Hd5dW9ikcAt5Af1WcFjX+RHgUgfNJN/tW385lb/tUN6F+2Kfvlm+rXoQ3XhSvtLjEzNyR0DO3b/jxeQL3+TA6BzVCvVuT1TPWl3Az12H8fe80XXmLnCze8T3jUWpZDXe4gM4sxeqwYOjwEWrueUK+RVFWP4jaA9ZJYbnHo5rM3DMrlHEM7Dp/bcYfcrWrP9i7v78ppbBZ2yzV7j9/lOobeeWjQWkCJvKLw0TkJXJo5AcCf1rdORGRgec4l55LnaZ5zzo/ioTu24sqY7MAPQAAicLbONtL1A3rlhee/9NSN566FF5+6+fTNI1bZRB7HqCa1lGmehzg4ot0A1FRBgJQISi2mhhCYfQmF1VId2u4Rb4fkoE/0ARqYgQCIc9FrMSJGHz+GZiAKvmYCsc0MphSZo5mpmIq5O40URVVNDAUZicMQNxXD+VwrRmVEwm9Pz9yJeVPS11cPetWqVatWrfr8azWgV61atWrVqs+3zOzeT1/PZx/DdHoxXYDpEDAxwvRQdg8G1oMhgQERhxBx3MAwQEigZlXKPJeSS8lqAgCBHLObp90+hbAdx80wxMDehWZIBoYcMQyQkqUEIZpUqXOep5JnKcVMqC0fV0aMgWKMxAwAyAEpGEdgMoaipZQ55zlfXJRpX+fCFIa4Obp2s1h4uMvvvP/xH/3p9/7+//R/vPXTex892Fmj5ZLJslR+yb4CAAC1IDQAEnrpmRFzjOnll1/6rd/6rb/6b/7V555/bhiGb33rW9/97nffevOtUisRjuMYQ3RUbpVacnGm82azySXXWjkEz5TO86SqiCRLPZq1LkFVzXluyALREFoi2MxE1GOeflh0yfEFkdY46Fb13FEeQ0rur/lRebA6cEjD4A4udF/NDKi5aWILgwJATRdD0j3GWotoBQAn/PbEq6+LdxCH5zcVEYk4peSFiuM4MrPb6NSq9pwiQh6ndRhIZzho/1IXh3G320/TVGvNOZeSa621VKk+2VHdtV8yzvAJ+xgfdQc/S/98BvQnX/rPZzpf1b9sA/oyBI6P+L9tKgPbFAh7d6GPC2Zm3IzbmBIRhS5EwsUOFvEBHGN0wAV0mzhwm73wsGvtbPRmbPdboEj1genp48VQ9hvNtxaIA7P0RQDErKp5nkXEAGKMLXpv3YDu11hETBXRKc1YaoHGwyGfTHLn2fciKn4PWqO3mD0SuzZVTUNq3Z49lt7D1LjcI58eYN2Cb6Dwnv/tQxGREEW1iorUGEOMKaVERCp6/8GD89OH+7MzxyWbXWFxPDIgL3fKjMRooqjABgHg5ohfegx/77VXXvvynWtjOt4OR5tkWmqZ87TfjuNmHIdhEFPRigHVpEo1ADA0Y0QGIL/WVcTT3CIqtSLhMAzDMMYQq4hoEZlVZZ7zbjfFmJhY1BCJQ9xstqo2z7NKNRMC6x84Boa+cMaMvLeSGJFBTVWl5mwYeTyi7bVZtZgBw8MHN0N6WOni6//Zf/crjP9Vq1atWrVq1V9erQb0qlWrVq1a9TnWu3/4jeHm84+/+rUf/5O/a5aHSIeB2UrdndbplFRioBg5phRSpJAErKrWUkVEq1Q3G1RCSjENwzCIl5KFEFIKMZAq+dp/aQvTkQiIlbCY5ipSs0jt5FaMRCmlGCOYISExUkgQGBBxnnWa52maa8kmwgRMGDkQhxBCGGk4qsofvvvh93/wxre/+4Mfv/3zN3/ywVvvfXSxm3MWBGiE0keJC11ueyN2wAUS3blz55Uvf/m133zt8Sce32w2D08enpycnJyc3Lt///T04e5iBwBmNue83W4Otgc5z9M07/fTwcFBCKHWWkpWs3Ec3XSrtZiZ010dtbEQOTpmF1W11uLWUill4fC6yeUU1J4WVU9JxxCgvVA8KfkJPHQIwWsCF47q0sIHgJ5l9X2FsDTO4ZUiNUR0NvQlVeCKi01LMhpg4VBz95rbavrOcm0Vee4GMlNKKedSSnaARq1SioOai59AZ+92ec2gY77dsV7StPCo07dc109d6qYrPIp/kQb0L9rdX+A5n2lAf+qFnz76z97hpzf1//lrPH7qrwjQJyUQEBeABwJzYA7c3WciCiGGELlBPKCKIEBKidmRyrCMfEIERHeiS60qombL40somoh9nsMd8GVAxBiJSESwTTCRo5y1Vz5KrWrmTyMiIAaD5QnQI/GiLVhrDeDh9Zt0Zdx5pBdSTO6M+yiTNjptsZWHNDBzd7m1B77BU9d4peGwXxro0y9tXsqz0qri6wmWzytTA0BqtZBmZj4XINKmY/a73X63m/d7U2lXHREITRW8ErNH/4ka4gMVGIAARoajhI8fHz735GNf/coLv/HyC6/cfvZ4wG2AiBIDBUYmMBMzBUJjNg6qWKvNWdAHALNPPIgKmCFglQoGIUbvwqxSVYpoEa1ggBiY2MxKrT4bNwwjgNVaVVRFpBYpVUWRMIYwxBTTgOB8cAREYPCYuQkYkFHA8aCanZw9fHDy8Pwsn8k+GLDq7/+tv/NL75JVq1atWrVq1V9arQb0qlWrVq1a9XnV23/8DasWAWcLTDWmsAEI9YLzac2T1BpC4sAYOQ2JQwCiXGvJuc6TqrinYYhGFMYxpiHFpGoGyMxGKAgoFRXICFVBVbUagCEgk5jWWkWllU05fJY5xRiY3Wg0ACMGIkSy3U73Oy1zVakIOo642YSDTeIQwxDi9qOH0zvvffyn3/rOn/3Z9/+fH/zwvffv3X+4m6RVbxGA+lp+AGg23oJFNScEuBt7eHh48+bNx5988s6dOy+88OILL7wAAGdnp2+++daHH354cnKCjRnhhAqbpmkch3Ec56Z8eHgYQvCmOzPbbDZm1nGxBr1OcBgGx0p0JKwtgWWvhpumyfEancbb7GPPfqqKk3k9/mzWgpPQmtnU/Vk37KBFLCWEQMTNURPp4F8qpQJYCNFBtz1/3SOV3URjpgWV4BiPbsCpl9flXIjQF+M7uLaUAoAeiL5iW2OtxY8553me8zxPtdZSqmfIS6kers+5LLyFdhimV2zYBUgCcJVDfXmV7Rf5z0sy+l+0Af1L9SumpD9tQH/WC3/FX8Y/Y4f0C3fb//Tc76ObaMjvy6JFfxSJPLfPjAAhxBATdVyMmSHRMAyBO+q9Y2XahEmf1WjJ+r4+oNdEGjEjkk9gdAPaAMyjzT6D5X1+BqA9zs+hRfWpY3CQAyytiX4WGhZGvCewQ5yVWgufAYCpllIAgBqKBP0ecQj1cjBmBgY+eySqXrPZOeyXpYIL4gMdSaGtofPKSEUwE1U/P9YPCQyRKIaofQqKiZzW7Sih/X6/3+1252e1ZKm11gJmQAtWZOnDNCRrKBoDNCAABvAY89Fm+I1Xbn/5znMv337m9mPbZ25sn7x2sEkUWEEyWEUzjhFjgpQAoxoVBUBGIr++fnf7u0cDIgoxIoCBiVYzAVD/+Ipx9PO2fDiEwL7uAQ1NTavUUlWECGPgEEIMDAZSKxABkiIAogJqNTNsDzLnOd87eXD/4dluFqgZdSAdDuz4r604jlWrVq1aterzqdWAXrVq1apVqz5/evcPv5EBAI0Yy2whwrWD7fEYLj7+ue4fHAwBgQCZ44gpQYrYUoFSaq21aC1kQEQpJRoGHDYQAgCgqBmI6O5it5v2U5kCcwBmoIiMAKKl1mpg43aMKYRGiPankINiQURrnhxrmmsrIFSQXAjk8GBMY4qbEY6O8PAIDg4hVytaKv6j//OP/8H//I//l//1j3/2wb2qWltUr9krhKAG8shp8EauFuRUNQBNKbz65a/8a7/3r/9b/86/bWbn52fvvvvuT3/67t27d50hMAyDW8/YURgewBSp0OESAK3QzFOTKaVSyjzPKUXnb3gy0Y1jt13cWfUzQoRmIFL3+32M0V/ufq5HI8FRzqopJTMTqTkXZt5sNgCgqqUU510Qse+i+3ROrTU/Nickd0fPo8rcbaBgHQltZqWUEEII7FnpUqp3zTGzwzEAIMYIgPM8u+VdSokxbDabec6eVJWGYmicjWma5nlyinPO2a93KUWlIiAyaa1mBvSIT9pswyv0lEtSxGIX2qcz7p/6lXU1oH+RAU2X/YSm2rO0n9jTpw4MG+MGEU0EiYmD9o4+tyDHcQwhBOY0DCmllJIPsBAuiS6+3Y76VkRUUyeSN6O5sziWg/SAsmew3c51x/nqtEStFRBbKSiASjOM25tBdBCNJ5evXn03romolOz3rEf1TS2lxIH7pAgg9XZNDkikKp5+dmpHCBHaoENVNTBmdgO6xbfdhScEn0BS85JGry7UNoOFTkDxtx9jdM61WruLCVFUdhcXu93F7uJif3EuJZtVQG6ndjGg0QCN/RNXu/vMZGpgFggT0TaF3/7Srd966Zmvvvz8raPNQQLNFyg5gG6PDigNGmIaDtPmYNgcFNFSRUX85lTVnMt+v98M45CGYdiomZjXioJnuImYOS4LI/xT1Eyd4R4wBApMDTiOYKJVpErJUquKcgzIpApzqVPO+30GpBAjk0OEEDjOuZ5OUxarYo/Lc/t4ojT/jb/5t3/p7bJq1apVq1at+sum1YBetWrVqlWrPmd6+5t/z6JE0nOAiDZEHJhIBct5RIkMkRkRAYk4QoiQIqiCia8pV1WpSohEzLHBH84uLmotQ4j/L3vv9mPJdaX5rcveO+KczCySdeGdRbJKIkWy1ZpW3y9jeB7aBgw0BtMD978wDwb8amP8oif/A4ZfBjDgNwPty3h6DDXk7mmO2x61mpJaVEstUizeb2IVybpl5jkRe++1lh9WROSpzCwySRUlahQfi4XMk3Ei9okTsfPUt7/1W4NPXQogcWBEIgCncBAzpeRoUs/0EhgOWT+r4vnXYqYGIKZFtKql1KS0aMIWECJjbDkwEAFQWJV6dW996aVXX3nlrdffuvLjS+9cevmdN96+sr/uvX2VAjjCYoKpGgyRWTBAYgAwVQBcLBYPPfzQxYsXL168cPdd94QYqsiNGzeuX79+9eqH6/U65+JWctu2Y74YpkZtntz0pmEiyjwgJsZS+kEh8JTYdX/MzSzmAABuKsFgpB6kjN2x8pzyVOw/7mFIQ7sx5+RZVc05N01KaWiWuF73wePlzL7xCBDA4tjoEMaAMzMTgPX9gJN2a15UJuSCG9eeA/WXMI3To4vO31D1sCqVUv3rIXXtb3Mtfd/XUkSH/0Q8Mare5A0QzYZGbbdev7eFakwo3pPeCZst3z5eJ9ztCVHLJ9vbMfTqo2b5yT6NH0PqOPJE3xWO/yNsYFg+agie6x+fBDaAJsgGBvGwThMCExISsgeJvX1h4BgjM48NDEMIPBIyzBPSIYaSSy55CBGPaxKmTl0een4S0lhLMNzofhv6eMaI8jBYEQUzJPJ7GT3d7KCYIfntwzePbKsqIhCSmqporTU1DYdQq+i4zgQIUmWCXI+p5gk742cXvagA/YwZ6EjSsGmAPlUdUE6cv6HerI+QREXNQmCfcLztpxvQZlZrMTVVyX3fd+uu63LfS50qMGD0oHW6AgiJhkasBma+NBcIz5xaPHR6+di9O088fO9j9959705qIUfLy0UAxgLATUvcGMYQE3EAVJFSazFAUzA1pkBAahBCoMCeUSZC9roWA1EFM2Lnepuo+m+CQCEQMw/sDjNVqY6YNlCfH9S0Vq0ipWpfhCikmAKjR9SzcAUWIkNUZEBjpV1Iu5reLVtfm6PQs2bNmjVr1i+UZgN61qxZs2bN+kXSj/7D/x4UYqW8rGS2jLiVCPo96fdr7XdOnWrbhdt/AABAiqhEpmLO3jUwQMRAREhkhFZr7bubN2/UWpZtC6ZmCgipadt26cAEVDVD4BCXS0NUM6tiVaAKqKpILUVVREqVYoQQAjArogK2i612capt7gJiJYCgZtVq6fZW77zz3ouXXn3u2z/83g9eevHlt27slS6DALj7DOheCkwOzuA8uQyJOcawaNut7e2zZ8994Ytf+OIXn3jsscf6vn/33Xd//OMfX79+fW9vr5TsZFvVwYDOOYtUM3AWrpNCYKyyF6kOnK21eje2oXifyMYuf27sOvLYabMw5jR9G1UxgxiDEzAABhJ0laqiAOYRbAA76KhmQ/dCACilNk3TNA0AuAHtAc8Qgwxe70Bz7vseAMiNLRpwHADQdWsA9E6MAACIUmX0xH0w7IsNYwycnQoCADB0WjNVGaKsomZqMjh3jnze2P6Qo/n5/Hj5qWPLn3ZXJ4023ybIfOiIJ0FF25HBH23haJtQjk8mPOKnD+DoGGOIjgmOKXpa3/P7iBhjWCyWTrdRUw8Lj8USwzXpRQMTmuWoAU3MMFJpYCDAVPOA/8bwEAYc8/hibbpnNzdTkVJKSA2HOLAjzFJKOLZJhIEfomCG6PucFo2mu+PgQMwh+urdxIw28DT0pnxBy8xE1WB81QOzHplGgLtBDIEDq2rf96vVul+vS9+LI9TNCSdOJPIakLE7qIwrdONSnQEsI5xp4alH7v/Sw+eeePDu+7fD6QVutYhkxQQCqVGt0Cy2mrYhtlpzydmQEIiAwUAFapXUtKlpFAxwmEPAQEQHEAoTgld+WK1SqhAiAcH4dg/dIM3D4YaMIlX95SAbkigQBeYYraK8xwAAIABJREFUyM1+3FuVIkBN2+zsQKRezCqA2rdX9z6a+q3c/MnsQc+aNWvWrFm/OPp8/gth1qxZs2bNmnVYrz37bA29YhYsjNBE3tmKVNd1//2GIMYQmoY8xQYAZqAGBjnnddeNwdWSSwWi5c4pN4lqKVKrSQ1MMXCKgRAIATkgEiEOCFQ1M1AkYMq15lJKrlLFRFHNPeitrcVikUJkTBFSAuYho8sNcUu0WO133bpTqGqSS3nzzbe//Z3vfeMvn337nb0rH672+lLVxEBHq2iMPQOMIUw3VA6C0Ahnzp790lNP/epXvnLxwoXUND95991XXn7lvffeW632x+AkxRjcY2IOTdO0bbter/xbxxY7g9Xjz7XWnEvTJC+T96NPQemcewBwV3rAAtwKjhhSlsTuRDvx2XuviWit1UORNNJynQ8QQhCppZS+z02TQog4cmZdCAiAplKlOh+DmVVNRNQGLu1Imsace1VdLpcimktGAOaQUur7vtQCBlOjOUcfNE3yM7Ber3PuVa2O8taCXdfXWlQVpnjqRkx1w4r9nH+q/KU0oD9j4dDL8CDs68sgMTp7Jrk73TTJV7xgww4eOBUwJIVrFanjWo6qk4hVxKP6uRRC5BCGF2pWShlD+t48j91WBgDfuT84cJLNPObsT/ciA+SAxGNeHHxvIQRCAgRTK7WoCIehTMFd9c3VJi9o8FAzEYcYAMDvfQDw/RzShBPBMZTtlvTBKQUAgIHGTSMhBCyXsr+3v16vS+7BFEwB1N3ncQoys43WnH44MEZYMJwK4b7t9MR9zW898/hXv/TYmbvaNiGSFsmqAkghRC+fMFA1NYVatfQFjQiZQoipDTGKqaN4vPgDAGKMxKRiBoBD9now1kutfd+bl4aMbS+BQE2rVkQIgZdts1gsU7NUYFUQNTRBAALKVXOWLldqI7Utxebmql9l0WDrD882W7uxyf/Ff/0/3LnLedasWbNmzZr1Gepz/k+FWbNmzZo1axYAwKVvfZ0EKbf94iaZpEiLyC0rWweWIwETMpOoekK21lqLiEjf5y73cQA2BwMj5sX2FiFYldz3ABaIAyHjlOtTGTN8XtSPRoaoAIIDmhmR3U4gh5/G2CxSioFB0NTASq2DgcuRuOW4rILrrnxw7dob7/zk5dfe/NGLr/34pVdeevnlmzdl1alM/bTw9t7eEO3D5WLrnnvuPv/oY+cfe/T8+fPL5RIQb9688f6V969cvrK7e7OUgkghuA0Wur4vOTdNG2NApK5bI2Lbtl3XlVLc4QKAoa9flZgiMYNBlWqqMQyEDbe3nAZrZjK6YxPQdjKg3Yx2DzoOtpSUUogHUqzHh71FYQisar5AQMyBOYQoUqsIAHh1v6eevVUaEcWU/O3KpSBiDIE5AIJ7cGbWtK2q1lLVNIbQtos+95uw2gkGIqPW63XX9VVqLYO7JFJFpBZvL2aj9X9IdvDefK51cgP6hHu7U3v61Ab0bRAcHz+OzwyQjQOehoaVFaYRzBFjDDExUwghhkDExBQ4jH07VVRVjKaYsXMwVIkIpi6F463q1y4AOCeHiTgEqTWXgqMBHWMMIeCIv6gikxPqBjRRQCIDm/bpLyKEwMSATrJW5mlt6SABrWoidaxdMESe8suHT8jGWfdMtINHbKLXA8hojg/uvCq4kz9y6h3pXnJerVar1f5qtV9LVqkwFjRMYJCpSmTsUGgEEMESwHbAs1v8xCNnn7pw/5MXHrp4/oFHHzrHVBkqWkVTH+I4VjYDqQpIiEzEjISE5vPkaECrWUrJkfTj+ocX4BAQKkAVR2kPuXJfVlTQKhXQmLCJIaWWY6NAIk5WUQJgwj7XUkXUBFQJebHTC169urvWUgQIDbvSrrp/8rX/+U5fx7NmzZo1a9asO6/P/78WZs2aNWvWrF92vfY3/1qNlCJjNsImpmg9y15iSk0MTTStJhVKLrkrOZdacy45l1ylVBHTre2d5db21tYWM3OgkNhKkb4rpRBRmxqTarXWUqXWWmufswIaMiITBqIATIpWTYyRQmjSIoToQdqQUlguFE2lQL+inC333Xq/1mpAwAlDotAqNjdX5UeX3vjW3/39N597/ocvvHntxh4zlmoiNnAiACas6ZQKdAtGVTlwjGm5tX3u3LlHHnnkq7/xG4+cP9+k9MYbb7z2+mvvvfeeu06IqGq1iLteIXLfdaWUxXKJAKWUWiszL7e2cs61lKnMfwJoDD0KiXLJIpI4iEgp1VkBIcSJwuzZYZHqnpmTN9yVNtO+z2PbQxKv+g+BiBDRS+lx6pymbmhXD1TGGJyWCgDe9q3UambuXANAapIfpes6RGxS4y3U3HEerC4DNXWXvG1bD2wSkSmISM7FK+L3dvdW61XfdZ13EazFHWebmrkd9p2P7w048Rk245yfJ50Y3HwHdSKg9KczoPFk8OhjM9F6gid+KuEQih4xEePihGeiU5NiTCk1KcWUvBxhKMWoFYaYvxIRh2Djoo4HgBHRLyxmBjNRHe8yxzEDMct4y7ime82fOAWT/e4rpTAHHPsBDudFtdbqzjURjbj2WygmfsTRedbRmyave/AKg0OO9vREr6UgolKLiHja2mAIU8NQXYHTUAHA4ewpxMBMhH3f7e3vXbt+vVuvS84ixTaw2ioD/3oDlmJoSmAJgAHQYKuFe+9Z/MavPvm7/+jp3/nKU6dPxWVS1jVKBhUBRkAEpMBEAZCRCJDMAFXRzHCw44eVK5UYExP5+M3GNUvAECOFCIHBDPynqjAAj5zFIWCKpgaoQFX9CMBgRMiMfZ9FNMRUaulLUSPjNld9/+beqiu96c7N/f2YMsY//pf/4x28imfNmjVr1qxZn4VmA3rWrFmzZs36/OrZZ589xd2CyoJFxdpl3FosmqBYVyAdIZda+r7runUtPaioVABgphBjCJE4cmAKgWNDzAhQ+lxLVism1bwxHXifLUMzGqjB0PUZOcSmDRw5JootxAAEqtncCDNEcJOWPIJ348bV/b1dqLlNsU2p1socU7sEDquuvPfBtUuvvf3DF17/1ndfev2d969c27251xVRZFYRU0NPznnTrw1NCFc1PXPmzKOPPf77v/8HDzzwABHd3N29duPGhx980OfsgWJ3RgCAkJljztlMQxxMn8DstgkRISEASq2OwgBnCHh3NaJaq5oxkTtBKcaSS9/3zsdgZo9CpxQ3cMnqEWkzY6aJ0eE5UABwC9vbtXls06EfbhV1XQ/gzGhzF4yY2E0lVVEZ+hOKeo8138nUvQ0JaykGEELybQDBVEVlikJOJlctte+zN2asta5Xq5LzwGc1NRGDoYXghgE90Tb8oyMi3vYz5OfVgP486yPQGZ/CN/9YEMcdN6A3Roi48cAGWcKv+CF/T96sMKbYNE2K0W9Q8hDxSJ3wxKx5Vz0ivwhDCGpWS/E0tIiY3pImdki0+9S2MYHc8vpVSynEkUNAPAg4O3bDaxS8qx4AECGATVUOvpjkxQ0wwkAAAJGnwLKvBpVcbjlHI5NHpzvLb17EUovPCSkmn3+8LeGQmDYLxE4gIhq6IZZa+667fuP6/t5e3+0jsjedPHL3DR0ZIwIBqBkRNJHO7mydP3fqCw/e9eRj9z9y36lzp2ITNDIyxSHnbEowdJsEIjPw3yliOo3cHJRtAAD+i8D5/aZDMh2JgHBgoJiZh79NAYE8y24qNfd96XNZZyUKKTVt8Aw6mRkhxtTknPs+iyBypKapRrurvNuVCmbCDCFgXPbb/2RGQs+aNWvWrFmfY80G9KxZs2bNmvU51Q+f/dOMixu2/XC63rBF4u1lYhSQ/Vo6kUrIpZSuz1ILIjATEpKbrzHEEGgMCQqAqlmtpVapYiZgBgjed8vMEImYOURGANUiSiHE1DARIQFyRVMTs2LuR4qaAhqEEJkIEW7euLba30OAdrFoFksw5NRys3zzrXdfvPTG937w8quvv/3K6+++9OpPbuz1WUFhSNrZ2OlrU1O2EQCWy+WpU6fOnD3zyPnzjz/++OOPXwTAq1c/vHzlyvsffHD16lUiCiE4gHWgygICUK3FzEJkJkbEKtXUpnr2XDIAgIFb0hx45NjigFM1daYqItRSSilNkyYANOIQVzSDOvBGbEpGIxIAiIg7VgDgHoxbbN5C0J/rR+z73sbspKqWkpmJmdwaE9UYokMJaiki6lxpTzQ74iD3vZmFkPxxABhzilrFuwYWqVXNaqlu6NRSRKSUrKLDOQMAM0SCofGjjT3rDsdvfzEN6M/t596Ptow/kQf90V72oS+O/emn0O26UN4WG4IDOINTTN63MHBgjjEE7ys4EJmZ5eB6NjCLKZkDNEb6zQhcxqlUAhC9ZaivCw0G9AD2IG9mWGslDkQ8mbzgcIwB0zH8BwCI4ICQIU89uqk4NCPFUop74L58RUzuZeecDYAOmhYqBx5ng4Od+MKS+7NN0zBxKcWp0qbmhBAcJyJiYuaUkjdBvXnz5t7e7v7ezerLTmrTEh56V1VTf4TQBi8fAAASwE6DZ7b4/P1nz9+78/C59sGzO+dO7+wslwwAtZrWgNTEBEjeeDY2bUhp7HKIXuQxxqB1atLI6POwqtkmthtGJIhINVNDY29FKbXUWqpWZaLAIQREHtYjvRwkStWSpVRBJk4Rm2VRXHW5EIoGaPDMzfu6net1e/VH/+Jf/RSX8axZs2bNmjXrM9Tn9oP4rFmzZs2a9UutF//2z7SK5hJiswh294KXRFBXuezv96v99bqUEjg6hLlt28VisdhahhCQyEzA1FTUpO+69f4q516kgipy4BBDjEiBiZvlwsvAuWkoJWgbW68tZwwBmYEZarGSLfer9X6fs6IZeSpWQBTVFu2ySW0IsZReVDhETgtuFoZROWSjf/Nn3/i//vz/+fO/+O56nd1IU0A1MEQbum8d9tfcJ5oihw888MCFixe/+tWvXrh44Z577rl06ZVLly69/PLLxIyDjWvTs1y1ynrdeRcyDwuXUlarFQB4fb0jj30DEYkxxhg9DW1mKTWIWEoOIRJi361VZSRzAB50/AM3o7uuM7DAYQj1qfpHrNGAxqnZoDf3c5969LACEU+H9rZpogpDulARkYjNgIhjjF3X5Zw3/d8Y42KxcCTr5NpPf6/X665b933nwGtVT1SrmXo0cjrrn/k1/XPWnWzQhyfY1YkIGeBojY83oE+4t9vv6uAuO44mfSKP+w4vLbhFSuSIaJ+Ytra2UtOEEEopiLhoW79ldOwimFIygNz3fl/dIgCAg06ZPuKJg+E3lweoB9sayReKnIwxrB6R+7RDRz8AcNiE2QD98PUqAOj73lss+jKPiiEiMTlUxMxyzghII+RafTZg8gWwaaEI3ClWzblv29Zfuyej+74HhBCCiroV62tdMcYmxRSDqHZdt7+3t79a9X0/NVo0VSZm5qrjnGCymXwnAAIIABHg9BadPxd+7ZkLz3zx0YfP3RVNJK/RtIlx2S5FTdXEjGPiFGlYdTMVqbXmUpw7v16vESBwaFJy97/Ugkht2xKNaHBERBzoUCUTDq0LmJhDSu22GpRSa84qxURqFTMgRMIARn3ulYAiKZFRNKRmcco4GgIT6LLu77U3++bdvPW1OQo9a9asWbNmff70H/0/NmbNmjVr1qxfML327LM1VGNRzmrYECzZuPa6dy2xECMEBkIg4pgQyQxpiMchEAAOxiWYgolUkVqZgJgxBAwROSIxGqABeZMuU28xZYi572spIUYFExFURRMwqTUDQmwaDIyIJrnmvvS5SQtGVjEKTLHh5TY1i6r0k3ev/PCFS9/6ux/83fMvvXjprXd+clVEzTGvHoSbgsZD90FABAT0DJ+nC++///5nnnnmC1/4wunTp2/u7u6v9vdXq73d/fV63XVdHR2cwRBRBQRPQ6ta7ovvJKVUqyeYy6FvU0oxRiLyzo3sng3zZOaGEImw9J1XlI8EV8qleFc0J7TmkokocHAGNCKI6MTZGEElbklX1cEa9jF78nyyzJjZTe5aq6OlmXnoaihSReJApx3aqTkyxcykeghS/bX1OTvtuuQstYpW75k2HnkineAvThfBn0Z4G2f2Uzqqd9SA/lhn3ADAjrGNjxvXwd/H7+f4Pf1cDGiAEX1DvraDSDEmv81UJISw3NpyYLQXByAiIaqZ1FpqNVVipjH47NQOh3V4A8/xYjeAodDBDWinRRMHHDoHOmqD/G1VG5ZpJtiQLzuNRA4vbtBS8tTP0wzAcMg+e64ZfEjD0T2APd11RASAIk6s9rz2gJ8molJKDJGZu65DwiY1OoKeJ5J7YGJCHhfhuq7ru67r+2697vse1CcfElMbQtACB28fTvcDgy0C3tXgfXdvP/bA6V976sGnv3j+4qMP7SzaFAh9Zik59z0GJg7IhH65qIqqr94h4tCSUc18GlI1MyQKzE4uAgQzUNNScim59B0SuAdNxEgBKCEyAJqK1qq1ipfbqDWxiZxyzkqGkUstqoqE7fZpDmmvW1/f3e9LFaFv7537Uvjgvro3dyacNWvWrFmzPm8KH7/JrFmzZs2aNetnpUvf+nqRHHPqY0VKi0hNYO5vWlkZVCPmGEOTiIkIITAAgqKKqZqKgJqhGegQNXbbNEUiJA6UIsZEHJEY1EANiczUBNDUitRapRZVERPvX0dEiAaOjGDiGHF0PJEUg1GISMFQMSVKrXJz7cb6vSvXnn/+H7753PN//Tfffe/K7s29XsY44S22nE325/ggIhps72yfOXPm9OnTjzzyyJe+9KXTp0+r6ntXLl++fPnqteuEFELc2toqtYrXfQMe4C8ImYMZMAUAYGb3dDw/GEJIKeWcPbfojzBzLqXk4oHpMdqMMEYjmRbohfDodjICYKXqLwEAUkxEyBxUyf0uRDWz6dAHFjkw0eBhmZmqeAbUzAB8z1OUG2slB6oQ8QBx7jSmGEPwxLSaIUIpZb3uRKpUX24oJee+73MutZYh7HwMxsF+QUznOzLI2xnQR/Wz54d87Kjwk7xZRzfDjS9uQ3+2kd18y0OfvTxqLAKqAoiApRR3a8EsBK61LBbLdrGIo4iIAJw845AHv208+DwZ0GGkdkwVAVXEmR7O9wjMyF4vMhA2BqKOGgMbmIr7qcbsMe2B/O75ZRFvTujD8XeHJpy0L6HFGN3LBgBEYiI1Xx00N6CZaQIog5mvfg2MbGYmtpFBMQWykWgwuM0MDIli9HW01LaLZc6rZrVerXIuw4LTcAJ8lkUY2drTQwawqlaq7a9u3tztq2nFBtP2I/fH0zvNVsMoXWBhJGbisHkfkRmqUUpNDMGh81Wk9FmkiupExG7bJsbkuXMxVSWpLBLAFMBwGBIJuNFPCAhGJgGIDVBFU0iJY63REDBSqUW1AgCHisRpaxHMrl672WH93e13015ehfh//Pf/1dyZcNasWbNmzfpc6RfiHx6zZs2aNWvWL4Ve/g/fUBJEyAiB6dTOkmqn3Y0FYwocAxMzooGIlK6WXrV41hmACYmJkNFhn0gHmF4z6Ev2SGCIKaQmxDRYCCkiAoiAVsl9v1qxd9kyNQRgjoslGNauQ0RFrGhipmqm6nm6nZ2d2CyAAxhI1fVa/u77L/z1N7/zV3/9tz9+7b0PbmZENIBqAoYA6MABs4kDcAAYHqvo7amnnvqDP/iDL3/5y9vb2x9++OGlS5feu3zZE95IRDiSLgA26tlt6KJnhkimVkUHwxjRq/gBwC0evNVrm2r2TXWIRjptuVYzY6K2SYjoLpWqmWmMyWv2fc++QxzJs6VkZ27EGGFwwXQcoSECM4/dCxURAdB3EmPMOXsukmio98cBU0CqvmcEAFUrxftPdqvVam9vPw+RZ/H8u/mr0o9Itt6O2/u50h3kZpzcgP547/WOJqDpJJudGMFxePe3PBMNQPFEQWY7iuq48wnoDSExEpvDMRyODgaoRMHRwIt2sbW13N7eTikBYtu2zOz3NfjCDuLE3JhQyzpa0AczgHN7wGejIXosVYgJDFQ1xOCFBQ44RrSpMAIAwrj84+tzRMxMAGgKoo6AR586Ykx+E8IwObBXSBChiJiBd0ocmB7ju0RIPLZLHVLDA34aTG1qc+gTyrBYxawiCJhiVNWu669du7a7e3N/f1ekmsrme7hR8eB/jMAIrEFIiE2g0zvhoXPLX3/6wq8+8ehTFx5i3WPrIkmbUgoRFIek+ci29iqNEYhvpRZfHHNeESD4ssEEyudBKFK0FilFRNVAMaqCCDAaEQZmTg1yUAETBQECIEIk73SIimhAaliqCre11qv7670s616KNeceef3M+Xef+k++d3tY/axZs2bNmjXrZ6r5d/KsWbNmzZr1udD3v/X1qJYsVC6LNm1vLVpSkxVIz2YIhIillFoylIwgTBYiIyGYh6DdsDBDGxpyEXlpu9s0agaIHAJxIA7e2s77a0kpNfcmdTBgVKuKEQFzVQBAAuQQKDBGDjFxiMjsBNW42AKgvsuvvPzKSy+9eunSmy++8u5Lr7775ls/uba7XgsgESCY6eBaDGhWQEMEsA0D+uzZsw8//PDTTz/10EMPnT59j6ru7e198MEHN27cWK1XE0TUU32qSoGJGBBVhhZhAF7i7ZgLTDECQM7ZPSl3SdxIMrMQAoygZbeqJzDrFEIspZpKjAOoRGTwuFNqJrS0iLgn5c61p5jdPp4c5+kTl+oAaZ3C1E7/2GB0CIARD63SPMPusUcVKbWu1+u+6/Kovu9zziUXUXGHfOI/A5zESp30OflMiB/57U+55196AxocB6HT14c33tjs6AZ2+JE76UcjIiDe2vDS4TyIQEjkwOUmJZ/E2rZxZ9M95SnB7TnogyKDEYY+yYE4AKA2nAgcQsF2y9cDCNoQbSTLu4UdxrWoA2cZAc2mw5mqARgR3+p+DitfjuxAAOIBrTNCemjw370Fq+r0osYnWgyBmAaGtU3nDRzlDyPep5TSdev1en+13s85S62mdmslxIEBjWAIFhF8ZW8R4NSCHjx998WHTz994cyXLj7wyH13bTfEJihiUtEMwZgYAERFVQAgcDBvdeulHMSmAgY09HgEb1YoY39UMzMVUDEVXzdUDGaoCog64EFSA8SlVDIK6KwVAzAxU0NFQmIDqqLAidslx7jXlWv7vQFk5T/+7/6n5/+3//T6Pzw24zhmzZo1a9asz4M+J//YmDVr1qxZs355ZWZX3rq0uvnhzb1rSWvbxnu2Fy0LlX1ABQQrKmpq0K/Xte+slhgwRW4WiZgRSavWUnPOBjrUgrsVShiYPSPs9dujCYxSpdSqUrWK1JL7HsDaRSNVai1VFEMgDus+A1JKTYghpBgXqW3blBoMAZENQyd07druu2++8zff+vbfPve9v3v+hSsfrvc6AABFqAgG7q/pEHEe3SW0wehBpNQ0d99998WLF59++ulf//VfZ+b3P7jy6iuvXr5yeW93N6XEIYiI+0G1ekMvjSkCYhWRIW8YEUFU+65XNSJumgQGq9UKEJiYQ3ADer1am1lqontGTpJl4iFBaY5YDTHFkkuphQ+srUExRmY2A5Hh0M6E9bL6GCMAqmrOGWBICHq7M1VRdVfLybdcay21hBAQcMxUujFdRWRq3pVzLrVKrTdv3tzf2+v7PpfsHQ1N9cC0O9pT8KTO5Wf9mfDk+z+RIfuZjeFEpiqeZG94on3hyd6gO2RA+6DtNiwOHHEfx7vwdvi7n8aAPva5BkDjib1dQt+ImEJII5QjpRRjMMAJj0PDTDPdrwAAviDkXHXn9vik6hUJxKyqiMhEpdapm58DfnxBz51WRPKpwHPQAMDsBjQ6gkPU5zrwsLMfzAxUjdn50eLQa0D0ogoHbyCiDutI5iUVPgAc0ERgqiFG5sEK36zkaJqGiErvMHqOMYnW3Per9X7Xrfu+r6XWWm0gQRugXxjTqTZGYAQAjGgJjQTOngqPPdj+/m9++amLj5zdiS1psII1k2lAYCIAVa1OvUdCURMBCjGEGEKUWkyViGopXn+j5s79wOBGMELgAW1EajSk7k29GIVTMsCcS0COHHH4jSFVTAwUiDgAsapyCByb5WIBabm7Lnu5VkBUOiW6QsgG/2z2oGfNmjVr1qyft2YDetasWbNmzfp56rVnn0333v3g0//oh9/88wZKu4iLQCz7mFeMVUREzBkMFAIjMgKDIpqq9Ln3/F2tXtlNHAIyoqMqyL0LM3dVTQ5UqqM7ShFiijEWEUBq2oV7BAjUtIt2sYSYkIkYgQAZyN0CU+izGVblV9788G+/88Ovf+OvXn/j8nuXr13bW5eqooPFpZsfNNxPMfA44RAwVEtNeuyxx//wD/+zixcvbu9sv/rqq2++9dZ7770HB6Fjc8jqGCgeDEpiUpH1ulMzBNioAa9g5i/fsRXe5ssjzx5dRKQQg9scpVZC4sCBg5rWUmJKAFByduOeRpYJ0gCbdgNr0BAzD0wsMpT/T0X6AICIIzdWNhjT4B/DVFVUaq0TNxYRSu5FBi+q1lpzXa3XOfe11lJyrcXjjOan5nircNOK/tjPe8eYiYdAJQBgx5mgx212XLT20GZ2uzHdGebGsSM9+bMPfXfkmXgik/y2r/HwkU7mUx/z2OEXdYyZffR82m0Ou7mlHfcmHn3KbYjSR5929ETc1t8+0Tmbbj2/ZWJyIzqlFBF5XMIZDGKPKTOjqtVavVsrEjmo5oDRzOymcC3FzeihmR4e0HUABh9ZVfu+911P4GYAmPDQAOCzAY5PJ6LppHrrxAnpw+xz19S9DwiHuoeD7YeuhreImRxAFEIgwgkk7VOfqsTAIrJer/b3V+v1upasKmCKzGCwiejBsRksw/AnMbaR7t5enrt78ci97ZPnzz16713JcsuwSAxSEJQJtre3U9uIaRUTxRBa4kjEJmImZtr3Xa2FOXAIIUbmSMSARABMFGNMMXEIQxIazMR/V1VkNABRNVGDzg+zAAAgAElEQVRQQ0QzERVvvSuqhmiIphY4pBgIsCqsiwnGdanrWglRKqw47lrznp792te+9nFX16xZs2bNmjXrs9JsQM+aNWvWrFk/N33nL/60De0W7OzxzcCwTLSIzHWfygq1RxMzVM/WEXEgdOwFmkftSilEyIFVAYk4BtCNbCMCANRaSskjY3QwoVXNQ2diyDGmplEADCG0rWMfkDjEJqUFMqvU2q+AFBAMDcFAVfr+8uWrr77xk+9+/43vfP/St7//o729vutrUdOxB6JtJkBHw5VG+xgR77rrroceeujRRx89f/78ww8/Aoh7+6u33nrz6tWr+/srGsvSvaR9KqafDGiAgcXhgeLNE4sIRORB6TFWPDk+Q+G8k0kmj5iIRgNImQMA1FpFBQBiYDOtVdQGf/kQqgAMQgghJNWhO+BgI42p6Qn34Q/y2MhRxJHNVmo1M184UJXcrYeVgiKllFJyzkU8+226YQ5+xAc53djmszagNx4/1hFHPDqM4xzVacAf+8hH69iRfkodM06Ew376CZ94nPSEmetjtjrsguNtxnrMMY/ZDDa2tNt70JuyI1/cZrtjDOhPnZ4+fK0SEzOHGEMIIQTH54TAiOTlCMzBPVkz9Val48EJp/US9EwyqJlXVBCzTy5ONNpoHOrcdiilDPyNkdIOvp4kAhs3+9SG1JfHnG7tBrRv6dts7tm7DDqRwxnWvj1Moe4DbP7ADEEnXajRGKYe+6MGMy05d96WtORuteq6tVd+DJUxjpoelyX86vYguvOctho6d1f4lcfv/5ULDz7xyH1n71puNYzSoxa0srO93S4aBVADQObQEgUAMq0qYqpViqmEEIgDEvvsSxRMzeFOIYTAYQCPjLOwSEUER5v4tOeUJNFK/muQUM0X8DQwRw4gUkvt+2xpuwCu+/W6y530XcnP1y+dx7e27eaffO1//bQX3qxZs2bNmjXrp9JsQM+aNWvWrFk/B5nZlbde3L165fr7l5s2hhCWkaL2lPejdoGMQVUKhUicShUDQ4Iq4jYss+f1OAQOgQgRmYBD6TotxQbH1gy07/tuvY5NDDFwYIcjEzFzII7IgWOKKSETxIBNAyagCsiGAYBBJO/vra5/4O4zIBhYFd1frb/3/Rf+6t8/9zffefX1d66tq2f6oIpW28g+TwhTRLeJg4eoEWOMFy9e/L3f+71f+7Vf29nZuXTp0kuXXn77nXdT8pr61Pe9mRJ5ZNi8A5iHHiefgoiapvFHvPEXgHvB7MzWWsXMPKLo3vBUWY+IpRRVddMKAPq+Ux28H9+mlGKmTZNEat/nnDMxtW3rL8u9D98tIYcQzcy3hMHU9qr/A6h013WTH62qPgCA0flWrbWWnPu+k1prlVJqrcXbEo4ndBNQcBID+mRh3Z/GgLZbXM6f2oA+/ORP/nlV76ABfUyQ+WQGNJzsNf4UBvSRU/pTGdC3bGZgYCcMOH88i+MzNaCHB3FI2RPxQItuUtu2i8UypTTe436j+d9CFJgOWpIiojpYY+jXGgdv2nkZOBjQtrEC5De13+DM7Pt3xPy0wYR3H83kYbkLEZwa7zR5d659nD5FAYCpiaqqTLUWMICtdTyLhoiBg0e5pVYcRzsGxA1HFraaqcqNa9evX7teci9SzASJ/UDDicRhzwML24yIAsGC7cID93zli4/85//4tx5/+N57tlLCitJZWW21MaWAiEhMHCgkb4YrUkzE1BCBCZlZDapq7osZMQXvSgjj+t+4SDBa0CZuQA/kDQAmNgAHoRBxir7gJ1WF/DeLqNZScumrKUeOzY29vfevf3BzXarVXiBSpUb+6X/zZ5/22ps1a9asWbNmfXrNBvSsWbNmzZr1s9alr3998fC5h778Gz/85v9passUtpoYpYd+lzQnApMitUqtFAKHKOatBWHo8MQxhBBiDE3DYCBVpUgtUgW8q5+Zmqq5t4WGoEPujohCiCm1S+KIFCCEAZiqFdAgIPQry2sTFQERqFVyLn3XKwLEENvF1Rs333rn8vf+/sXn//6VH/zgjfev7++tS7XB/TIzcX9r09FCcGcBDBHgwQcevHDhwqOPPvrwww/ff//9ly9ffv/9969fv77u+jwYskPA0O0Pd45yLohAxG3bqsp63TnRYmdnx8PLOWe3j1OKni7MOZtBSgkAxuAzjBnDA1KEx6Wd8TrZQ3AQZrQYg1vDvuUAafZX5AlKA2dieJJx6kbo9fhTEDKEUMbqfne5zayUWkrp+77ruvV6lXPp+261tzfZVaqOSzlWH/1B7oRMA7iNAX3YuT7OM0QEPORx38b8PQwjPmZXt3viJ6NCGzgJ/ZjHN765nQE6DXLk1xxjdw4rFB9lu34C3sexh7hlC9/jsdvcakAf0xzxdgM5ROE44lNv5IQ/UgajP/gxmx3z2KfzoG/vd6PfaN5LD0J0Izp6Pnq5WLRt2zSNO8WlFOaISJ6JRsQ4mL8mIoAYQvCJtA43rF+EUyjZplCzR6G9rGFKQAMM1OmNeYa8eyGM889QwnKrAQ0AOYtPNeNJGmeaya5lAgMvhiAiJvYxeZoZcbK40aHPZkaBQwgppX7drfb3u65br/ZXq/0pOj2ew2GqoYFZr/7KI9lWk07vLC7cd/czFx/68pPnH3vg9D1bIUFesJKWvt8jBMdEMTNzwGFyAEJC70+o6nMsUYqpLUVqqZuB8elcqamaciBij2IPhSOeYSc/1VUA1Odf9PtVUcVqVUMyChSiIPalv7Ha388iFW27amVD+ON/+a8/1bU3a9asWbNmzfr0mg3oWbNmzZo162eq73/jG4ylqdRtrwyhiWE7xhb6UHa1ZjQJiI6G8DJw5gCEyIiBDD2+nJiYmTEEq1Vzr1Kk5NL3A8Z0LKg2QI4hplRFDQGYKaYQm9gsENgADUlUasloFUGITNa72u1brVKtVqvVjENIbQXaz+WDm7svXHr9Bz965e//4dXX3rjy3uVdMVDA8XCgUy33pmeIgAgxpp3tnfMPn7948eLjjz++WCwQMef8xhtvfPDBB7VWJAJ02EWdumwREQCamergE6WURBzAasxhsVh40DjnIXiYUlLVrusAgAhjjCP3GY+gWoeUHzNPCGkPVvvjtVYATSkBmIh6i7PBJx2gIoPlZwamBx6qfzEml9H3ycw6Ngz0ZQJV7fu8Xq+7rluv1/v7+7WWknO3Xk+d0zbM0mPzrXdKxyagb03F2lFHeyrW39js2EHZEYvziJCObnA4Xn0C2Xg9Hnl848GPNKCH/DvghjF366DwuLDxrZuceLgn9HlPEJRGPPxenHi3Rw3okw3s+FN9u6Mc/cmn8KCP29tgURqAs4XBVIkD8cBqYOJF27aLxWLRptQ4n4c5eBfQwYCOkYjAzDvmsSM4VMUUNhAck6abfaxj8HUJU7UJ0rNJ45n8aO/aZwa1FhgZHW58e/y5Vp+s0OEYBtORwXPNzOw0DsQBRr9xdpyYj0MPAFUwNTOOIcSYUgI1qTXn3HVd1+33OZdSpIw1Frca0MNjZl4AExC2Azz24JknLzz45COnH73/1IOnt85spYZrt3sVrDJ4I0f2KDciIyIjI6CKqlQ/nYCEFGVKQBMBQMnFzLzlooGpKQX2H01Wu5eYDFHoWgEMwcaUN5iSGqlCiImIFdTQIKSscr2rvQYIrEFYAkn4o6/9L5/82ps1a9asWbNmfXrNBvSsWbNmzZr1s9Pz3/xTLBG6JTb7EHSR4lZAW11L2rcMXm2tUt3NiDEiECKFxCGFkAIG8tZNpqBVS8kl9zVnRFSppe9TYA7sHawQ0RBjE5u2BQBghhggNsABjKCqVhWVddft7+0RGTNEgrLeLd0+VFFFMywCy527ztz/UDV6/Z33/uLf/7//7q+/89z3XtpdWRYniOLoQqGBKYyO3YYBjQhIeOrUXV/4whP/5T//5xcevxBjfO6551544YXXXnvt1KlTbdsCQKlSRUNgTwSn1MQYmIM7RO4y11qnTHHTJGZ2S8d/NBSkh5Bz3tvbWy6XMYaR+mo4ZvMAwLd3dwgAUkpN04TAItL32WveY4xd14nKcrkkQlN1oAcSqrrTfuBUMgXm4P0JmXkkOJcQOIRQq5OmwcvMAaDWIfi8Wq1Wq1Xf933fd10PQ97ZNszEj8iifoYf5I5DcPgwbllbONqP7zjewolM5GMMaPukjuq0Lz1iU95JA/pEDOiTjXQ2oD+hjuzNg7Z6KNNtSASbKX5VYo4pte2iaZoQghvQ5tR7t5gRp5lh9IuVmHHEaMBYSzEeGX0zr2PwZoQAMLYBPADBO4x+IGkQuj87Iel9e5+pAACR3UCeyDw4ADUOeNK+ChI4OCKZiBBQVByXrGZE6M1eh0lkbJsaQ4ghDKcN7YMPPrx582a/Xg9v9waCY8KDmJnWSr7WZBAQW4ZHzuAzj5/7na88+eRjD9x7V9Pvfqh530pPYEzITADk5RFOREIDEamllFL7Pnd9QaQQYtu0Tdsy83q9tnGZcKzaAQVQsyp1TI6bylBBEoh80XMIihuIkRmB0WKxCIGrFpFcpK4r8s49kNpeo5mBkO2ALLWc0T/5kxkJPWvWrFmzZv2MNBvQs2bNmjVr1s9Crz37bMa+Ul9CT4oLhiaFCAZ5X/I+gwYawnqIyIGZmZGIGYjRBE1gau+naAYi2vdlTJAxGKopETIjMYfAzASElAKnBFJAK5gBkxlIX1RM1YpaX+o6Z0Mi5pQSM7DzNImBgqY2F13vrp777t9/+7s//PbzL77+1pXLV29kATEAgEARAIpU8CQseaH4AQNhsVjc/8D9zzzzK489+th9993XpnZ/b//qtavXr1/f3d3d398PPlYksQF4CgCIlFJyU0ZVESGl5KbtFAgMgccUIY6UVXEeq4j0fb9cLmOMAOb9t9xPYfYYnfOXxQyY2Z1uVVFRHZPONpK0iVHNcaNiBuO7NKA8AIGZwXBky6qHGcd+hk7rJodp+EsopfR91/e92zG1Vh+5iIyWnH2WH9KOQzl/gsMdcpyP+NRHd4V4aP/H+47HjutTyt00O/zILd99NIYCb/mp3fqTyYA+yIlPWx460Mb+b/tqPvZlHhoqwIDavnXwh0PrtxnSMXv+1Of5mNWGo48cs9FB17uD5x3a7BiY+LD/2yWgbx3D4faYNmCKOTARErXtIjWtz7W+LuWMeVE1MxodW29CCABuTG8eZgovu6YCi+k1jpUQMiE7fIFqetx3uPks3/EwJQ4LXUOqmQaXHNxlBoDNug1fD5xAFoPZ7YANH7a3TNxAefjc2HVd7vuchz8O/PEENI6gIT+VaAZgaMAIOw2cu6t95Ozdf/CbT/7qkw/df1ebsGLtoGZUYYRai7/wEAIHRqJaq1SJMQUKhNF0sLlDDERUizBzSgmJVDXXYgBiVmrR8UUxc+DQ59453V7tU0sGNQRkikxMQztJq1JESxHpxWh5ClJbBLsiVU2q7j9R7rna3IPL3/gX/+q4y2zWrFmzZs2adYcVft4DmDVr1qxZs/7j17e+9fXd0u3UNkPPQotEyya0li2vVHtkIArIgTg4X5iZ2P0PZiDUrCAGWk0EVLwJloipKCAhBcLgmTokQEYmZkImMFQDrCJWC5QMUgHMVGpfTM0AFQgRUyAFxhipWcSmSbGJMREHRbrR17fee/fF7//wL5/9m+9890dvvP1hV1QAdbAiQN35BYDJBh7MIFwuF3ffffeDDz544cKFZ5758pkzpxHw9Vdff+utt6+8f2XRLkIIy8WWl1d7mHosjeeUopu2nn1218aDfiFEABMRRJrsmzFySIiOT0Vm8pwjDP7bEH92YHStgoiqAoAh8Ah4RUQMzDFGAKi1esxQQUXFM4duSg/7Gd9fIlI1E0/dmpNe3ceZvCER6bq+69Zd53HnPudsIna8z/ZZRwSOg12c9Ikfu+VRDvFh7/WwYXhbfYqE7OZzb//04UpVAABnInzMoTe+RYSh693mrkZTG0fD9xA45fjThnDYnD/2pUxbHDjOiEdXKY6+O2ZHtzr8lEPP+IjRHh3YcZsexpPgce/DEeTLMSPD23jQJ9uZHf6BmUkVqQOjWdVENYSYYowxojc8Hd3hYVZh0pE84wgIn6MmP9Qf9B0e6jcIYxmBA4XCkDse9uPTyCFHG4ZZdBgGqeeAnf7v0xr7DhV109QeDjfWEByk1z3NT9POwdfYpsMxh7ZdBA4cnFjixvFBk8MxGY3gl6EhoInhtc72c3fl6nthuV0p/soXHnjw9Pbpu++JVkkLSJWaRYqBDpYwk6iJWQqpiW0TWgc4TzefijGHwYA2LbUCooBzkIb30xvv5r53crQTT0rOaEaIAUNgDhxEikhVFTERk2qmyMaBF9tF7PreXpdz80q8+/Ty+o2b//Zrf/RHX/u3H3+NzZo1a9asWbN+Os0J6FmzZs2aNeuz1Q/+8t/khCWFppZAttVQsJLqeslAXsBOyCnGJgEHU5Ba+74rpQAMFdel6wJoGwhUHdEgombAMQGyATEnjimkCExAzhPNWnLOvUgxU5FqWkHFQBGBhopzjilR09JiARghNrhYIhACAQXD0HXlue98/6+e/f++/vX/+/KHq+u7uVYRQwUwN6BtIEVsJCwHGgcSXbx48bd/+7d+53d+9+zZs5cvX37xxRdff+31/b3VaDEnQhIVRFTRUooBAA1130SYc0akxWIBAKriUWFV29paAkDf5zH6J55shtHthcHlQeYAALVWf7UhMBETeVRZ3IN2y9yzjUNwTrVJDREN9exmHHmAtKo4n9pXB2B0oBwMohuujf9dq/g72Pf97u7ujRs3VquVN0uc+goO/s6xqIfPSseYyCdLQJ+IpGFHoBxHAtC+2Wepj0VDDG0E5cjjPNqXfiUTHM3qAgARAG4suYA/xQBg6hg5RFcnK/A2Z2+8lj5ShnDEqRz9zVu2uuXkmw0O7klP9nHYDfuoAPUxcBU72i/xKDDbOTMfvQ0cH4I+EY3kJHImPBKHGJumadu2bdsmJQBwko9XoZRahuwwYggcY/S5SERSSjFGnxOGCWQ0oCe8BgC4WzqtqB1EkodTMchnG0RiDkMFxmhkuyPsPB9EPJrFHsbMYSjD8AIM07Fv6mBSiyjY4UD6NF+ZqUjpuvV6vZZaEcBpQhPCaDoUIAAYmzHATpMePrf91afv/8e/+eXf/spT504tGxTNKwZhNA6oJatUQKAQgXi1WpsYQ3A2NAydG2spVURMB/ZHiAEI0X8dDIFxLbXkUkIY+vDWUkSEkBgRAbVURIwcxPHSaIbj1UgExEapYlit1+9/eG23W2epkjumEFP4w/92ZnHMmjVr1qxZn61mA3rWrFmzZs36DPX8v/tTAGYLpdUmxZ1Fu4gWpA9SgimYAggRApmBqQ0Wap9zrUJEIUbmKKUwWGJiRPSmSyJmyhyMyJBoaLYFJlWkSC3qQAdnFSMCoLsOhkDMTbv0tDUH8pJlN4SKAQCrUVfhjbevvPDj17/5ree/9/wL//DjS6WACCh4y0FUnOKFU9jQZU3b3nPP3b/y5S8/8cQTjz32OBHu7e29/fY7P/nJu1c/vKo6mN8iCmBEFGMkQoeoikoIERG8Ox8zb21tOU01594MfHtVzTkzD/XvIQwsV3/FKaWxXdVBhTszEbHbhTqa+D4SN3RKKZMBHTh4lnBoBRnJkbiTm6emYECEZqZmUqs5fwQARltQRNbrzs2prlt363XX9aUWERmzmRux1p+l/3xSA/qYR46CoQ/pNmwN3PgS4bYmIh3lTh98dSTQeuyRhmd9TI9AmEy02/586rh4rDfvbvKxJ2Oyaz3cvmFAH2s/nywBfQxZY3iptyV+DPv/hFfWcZcibvz0lm1vZ6kfHhIesbCPQXCcaHR2Bw1oAABAQCfzcIwhxhRT8phtDCGEQEyyYQSHEJwFJGOjQp9qaq2l1AnBMYGbJ3MZRpzFZgJ6BPbYsBoyoTOARG2cuxCRJo96XEIbOMiHXgvCwUQ1zlfms5/vX0Tx6G12kHMGBK1aS8nduqulDC8dDA8VLSB4W0IEYIPtNjx4bvuJ8/8/e+/2ZMl1nfmty947z6nqC4AmiQsJEABJEHfSIhWmTI88jHFQYSkcsqgYRvif8JvD4bEf+GRH+NFvfvHDTDg8hkIzskaChgpR0IWiKJICSQAEiQtJALygceludHXVOZm591rLD2tnnnPqnO6uboCUHMoPZHdVVubOndfT9e1v/9adD91754P33HbXrfNb5pywNGzzRAGBwIoUDBFDXC46yQUUQmAmRqJ6JhxxpF56l5iDISARhzCMgmAppe97vzoxhiJiaoEjGKioKXjcXv0+IQD28R0UkZyLISlwBuqlXFksFh2IlDSjLAAIv/mvJg960qRJkyZN+gVqMqAnTZo0adKkX5Se/srvIyiCCXMzb07vN/OAcy4REFWlLyYZQAKBSN/1Sx2CckXVACiE1MxDnJkomjFYCEwO5ZACKgAAhEZoqiACkq1bSt/2uXegBXAADhgScgAOwGyAFNPe6bPEwcDMMkhvuQcpJfdt2/YFjtpy/sKVv3v6+b/8m29/55kfvfH25d6QwRBgoFCjrsJwaFADvMw8m89vv/32+z/ykc997nO3335HzuW555595ZVXLl28pKoVlwwmosvlEobqf8xUivR9l3MOITgruZQSQtjbqwa0G8T+UxERKSFEN1aYAxG65W5m8/ncU8l934uI0zkQvS4WaHV23HLxoDTnnPs+AwABotcZQxh9IqMKd+ZqVbEnEJnJ++m5RTfBR2sp57I4Olq2bdt1uWtrPtrdRvslO87HdEIDeleQ+QTaQfzdaGMwoLe6sKuG3obbOMbGr9461St7op7uih6bHE/m7vaNT/ZPaFsNW+wosXjiphAQbQ0uvO472/rNtBYrHh3Fret4Mq1YH2s9XD//J4rDe09wK2m+K2p9wn5tl5d8N0JAHGEdREwhxhhCCM7lCDFQIJ8w4Rnn1KSad0YaiwFKUTegxwQ01MhzrRAIwyEzs7M4xmqHZrCqLeibC/j0C0RaXz/nvoKdEZwXMt6cNgSYEdGj3TBiMxDGDqiqlxrYPKWm5g6vIaEPwy0WC2dDl1zUMRlmq3Q/Vvd5/X9zhHN74ZMfO/fwPece+OBtZ+d0usF9hr2GA2HOPVCAEEtWHx/lUPn4GxB1Q2IPbZOCgce6VVSVmFW15EKExByYVdUMQ4giJkUQgxqKaB03YkQGZCSkvuvaZQv+4QUU908D08GibRUFKAQAIzb8jf/53753t9akSZMmTZo0aUOTAT1p0qRJkyb9QvTdv3xCFU0JyeKM9uezeaQAPUjWPksuJQsjRsYYwTTn3CEAE8cYQowcIhBTmmFMJoI5Q+4xEAKaatd3pRRmUpMiueSsJZuUgBYIiTDEhmNjSBgixgZTAyFCSOYTzzlYydq1uT0qXSu5d6itALz6s/Pfe+FHT3316R/86PxP3zi8fLDsi4B74lo9Q8O1IoOEYGCqAHjLLbc8+vjjv/Zr/9kjjzz25ptv/PCHP3rhhRdCYDDIOYsU0RobdMeZiJqmEZGcc869wzfMQKSUIjHGlKLnnUWkFHG3ou97J7HOZrMQgpmNM+JjjE3TjN863NmdGQBIqYEaaq6YDhE1sxDYiczBq2URdV2nqiEEN0dyyVZht/W/PNTX8rJgSKSipWjfd23bLpfLruv6vpNSKrK7GpGKRG54VfTzTdtw70r/xA3oayMvdAWd2OBrHN/TtXsybjg6rTuIGX5sJ0BwoMGGAb0dKK5naWXODusQ3pgBPRTB3H1nbp//E9jQ77EB/d6GoNez+e6EIpEzIELTNHt7s1On90MINqCcmbnt2pKLz71gZvGYsNoxA3ocLRsdZOZKAVoHbtDxkQkcb0BVJaYQgqmJqkipZGpAf6s4rQhqPUPzewyduYxE6IOGK+JHpXFsXrJqfJupqZnPC8Ehk6xvvvHmwZUrbm9DzRgDrk1I8FeaR6EbxHN78eMfOvOpB9/36Yc/+sFzp6A9wH5J0jNhMSgGMTZ+zKqlBqyra45gBuoFcZmZRQogzmZz8dFEVUBAp+KYAUDfZymKlVgC6nAo8tiznwqoV9Uz6b4rIgtRuLm8bAtGC01MISrIKetn1t9mX/ziFIWeNGnSpEmT3ntNRQgnTZo0adKk91hmdv7V5xfvvHl4+S0DaSJGJlke5FYKiGqxIqZGyBQCR6ZIiMxNwhrYwuC5MAPNveZeS4GSsRQBT+ZyyaWIQmQxK6JIzInAUozOmqAQGw6NMSMxEgOSAVjfqUgRKaogYiWXfmlqiKTGl68sXv3Z63//7Avf+u4L337upbcuLRY9iA5Tx9diljZYc86dCCnMmtmHP/zhj370Yw89/PD7zr3/4PLl1179yes/f/3oaLG/tzc4uYGMBnOBUgJmCiF60jmlNBrTjs6YzWbMJKKIwszzOQNU4IZPY48xOj3DJ7Y7ntWRrETIHD0ibVaNy8BBVU0VkWGoMwZmZhpDYCLwIlfMqkHVmMnR0mo+Cb0eu5kRktt6nkbMOXdd3y7bruvatm3bZc59KQXGAnBrQUUcT+IvJAV9Eo94p/v83oQSNmzlXb7qWrB2dwPX+Nbr7q0t3wnsWLfXjvMorrHjzX6tGrGNLU7ewtjn2lVcj3keW3eLmXxsF8dPCo73Tx0RcV/fVsagDT29DuDj2G24+nYD+XGNi3aC2wZhVwp7l4l8kgcC39vnZnVoBoYOQTIHKQuYmBUziSmFEEKIjukIzEXEVJkDMxURlYr0QYRaqhQgMKuZqfpbwgf/EOqlMl5xL4ZjGlgYhOSbWI1GAxkDEgVHl3jRVVsbwSIixHFca2jTDKna2QPfA3RVcXM1NEJYr4e/sQyQORAxouzt7yMRALTLRbdcqunqo6A6xu7bgxqIWr7Sw/krwmBx/6B93523zM40PAs2b7iodkWRKBBFDlBvAh8sJnEAACAASURBVGRmRFIVb84QiCgyd12vaik1pRTj3nImopiiiaiIFo0YQzIiryKLUhQAkZhCIEKrM03UzBCMAJnQzIoUYy6gMgs8P00xZjUtRZfa36Wzt8uT//t/9Zv/3Z+8hzfZpEmTJk2aNAmmBPSkSZMmTZr03upb3/o/zp1+6N4H/tl3/ur3E+gsxQCl7w7z8ohREA0JCCnEON+bN02TYmRmioFiAEMTga5HFRCBXErf5b7LuQdTQuhzD0SzvT01VCCKUZGMqJk1IUVipohAqGqIgTgaMxiACPS9dUtdLNqu7XK3zJmYOQYzC3HWzE4tO3jxhz/58lf+6qm/eeaZH7zWG8imRTTYZ6hgVv0ONIOQ0pkzZz7wgQ98/vOf//Snf/Xs2bPPfOeZb/zdNy5fvsIhnD5zppRSSu771ieGxya4FcdD8M9LgblT7KgNJ5w2TTKzo6MFADDz3t6eF6qKMfrcdgAopbRti2tTzs2g6zoAaJrkMcBhYrtVuGnuiQgBDYyZAKzrOp/nPmarV6lVRDPLRXS9zKJ5VTFz5kbO+fLld46uHC6OFn3fFykieeu+wK0vfhE6YbR5x4aI18/JXjPafHyv1e66WoAYdhWmoxNldQ0H3+06weHN6nlX7wwM9vB1Y7knyYDvXGcdlXC8l1tLdrawY0OtUJdaZY5Qxa57CNdo+SrbXrMI4fVbv+pej48u7FpzV5duNv58sqZ2nHzCGONsNr/llltOnzo139sbiRZ+5p0gn3NWdY4HVr7P0Ja/0IhItXrBXsV0oAlJfUNZnS2BREOKuYZ3Rzx0ztnMUmpCCIjUd72qIlUuhzfoo3SOqmdiGFj2BgZQX4gAMBbqXD9kM3NgPiKaSinZIUVEfPHtC5cuXSwl1xkkBAArJgcgOJRDASLCnOG+O5pPfuzO/+LTj3zszls/dG7/7H5Q0L6U5XJJgPOUUpyFkCiEGBMid/3S1AigiBBiZF4s2txnRCqiWUruMzM1sySlSC6SCxExcQjsByBi4HUCmoaZxBPWKqKCZoQYI5dSFosjigGYi0KYz+P8VBZ56+Kldw5zEYFTh9pGMfjt/+EPb+Y2mzRp0qRJkyZdRZMBPWnSpEmTJr1n+trXnohYMF5JR7cDlMQYLAfrGQqhhUAhUEwBiYgDp0hMBKhSSi4l577vpc9aSqIQCFENTEDFTBCACIiYY6DYALMRY0wWIoRITMiEzJZblV7MCBkNuz6Xvte+JxUsBSS79dqrYggcmxBnbYbLB8s//crffO0bzz3/0k9ff/udi1cWvYHa7rChGyvM7FbFpz79q5/45CcfffSRw8OjixcvvvHGG5cuXjo8OEJEYibmUgTQYgx935eSOXKIMYQgOetQJNAnYbutU0pRFTOLMTqRY9yzU55DYCJGxK5rc84i0jRNSgkAuq7vuo4IQ4hNk/wAPBJqaqUUBCAc/GWs8AOvJwZrRs+69SOiWWRAtVIIzBzyoKOjo6PDw65rS85OiXUTaVeO9Jfwj65/FAZ0Lam2ga/AocwaVM/rpgzoahNf3YAefTr/buPuvaZ3/J4Y0NfY/Bob3jSMYjzYwVHEtWJyN9nazp+8W1DMblv7H6kBfVzouWViophSSqmZzebzedMk5mBDfUJV9cffLeW6KVYkhpm5jasKpitvWlX9+tVahEOJQg4BsEKi3eYez8YIkmYKgJT7voioSoyJiETEN0kpmpnXO8Wh1KoNMzBWD8hw0tcHSCp/WQUMCBFQiTildHjlyuGVK13bioqZrj3Rq3OFAEZIAGx2Zka3n5nfc+7Mpx+641cevuvRB+49NU8AYqXX3GvfEzBx4NSomhQVLYGDf1KYWkDqezG1GCIGBiK1yrMWES1FcyGiwMTMI2YDAYlIQWHF4ak1Gb2vDq1SrNFoCpFizMDLvrt0+WjRqYiVmDFHLOm//tL/fcO32aRJkyZNmjTpKpoQHJMmTZo0adJ7o2f++o+y5I5hf3k7EDRNE02wLGaEMTQcmAhDoBhD5QGLFCnqod++y11XcpEiJgqxgRAJAYkd+UmMFDimSMQACMzAbIaGoKomRcwKqOUOtBhVuES7WOau11xSCIGQGDlFDkSmwBEoLTr70WtvfOeZl/7jU3/3nedefvty75hPn2V9tcnuzHzq1Klz587dfscdn/70r957733z2fyVH7/y0ksvvf76eRWNIaUmoap0XZ97BGhmTc45l8yFuO/dRDA1T+2pqoq6S+KM5pGvOkStzaN/dT4/ISL1fa8qDmz1XGHf933fxxgQsW3deK6sVVMtOTNzSklFDcwtIACHQdccom8yWnrVWtKaaHR/B6Br27brur7rDo8OF4ulSRn6djVYwS/IfT5hs8dW27qqN9C7ExjanjXedsIBKrVlNz9jOH3Xbt9/egybu3HW1+zvYzCM6/X8hJDrY2a2wxMqmGYzc3399mwNwLDqrm0ssPG4Nh3beoB+ow5/3NyNZoMFv9Ez//tkQxhb2611dFfJTTw+oLG9HzNbO9N27O9fokxVVCWX3LZLXhzt7c1ns1lKjb8nmLleIaxur783RGS8CVTRWfT+psIhAU2IXluv1i1ENEQ1BRtejA4vxoqNJiKvsCqoiCyrDHUhooptNmUhMyul+Ngek1dMHC6xx5YRjkG9/S7yOL3kDOZfA5I4Lj/GaGAl5yJlcMM3rodhZXGowuWldt3RhQtHXemOcs7Y3HnbqdMznLOxZu1aLQqAFJMP8PlEGGYW8XoDqMUAUGLhGDGEWifRTEVURUUDkQghFUIkQD+xzNz3nYigW+lEMGTDVRXQiElUxNTUSBRz7vpeQhMZzbJC4JysxNvuO//9v3z0wV9/7qRvhUmTJk2aNGnSNTV9ok6aNGnSpEnvgZ7+yu8jE3MUkTCjWROoLPYi7c1iJPQJ26IFTBEs913uu77rRYqKAAqogGmIiZDNYJbmMTbgZgMxMnATeW+GBCACbQfMZmBHi9J1OWcr0vX9ol1QDNyElCIFNNRlu1QxhHDq9Jlm1hCx++BqChTbHr/3wk/++E+/+n/9P3906TAvWh0dhQIAg+O1bfjM5/N77rnns5/97Oc+97kY049//MpX/uwrFy9dLKWcPnVa1XIuSAiAarpYLnPOXM0FokA+Yz2mGGNMMalpKaVtOwQgWAVRmcmzgUQMADn3zCGE4BE/d0NiDCmlkd2BiCEEZlKthvVK6wa0qjtuqmKgzOxx5tHvliGa7XPPFYCYmTjnvFwuDw8PF4tF17VS8gqNbau49dVt6PdW12JKrK11ncp+vtJJEtCe6NQT2bh4jbj0zqwruPt2gpw14vHGT0ixOLG/fDMakvarnhARbhnl10Bw7OgeAgJeDZFxDazHjWrwsteaWm/0htrfse6uDPWNdXnVAg7Qh5s86o2trpWAXp1ePFZ6EYkwhNDMZnvz+d7eXtPMiHm0ekMIOee+zzn3vjczBXBjehPB4fANIp8LYgDO0tChA+4pl1LGyRlOwO/73lHHRKSmpdTBM393gVkIYag9iO7YIqGDhupx+19oUOd5yHB6qm1bcicipuqb5ArWJ0Tou27ZtqUUFYH1uqC49qcBIQSERNAgvv/M/Fcevv1jd56599zeHafTLXPei9R3bSnZDDnEGFJqmiLa5xxTQxRUQUXBgDkQkSEW87Pg4wHmXrkzRgiRicDAR2zb5bKIDLUMGQhLyX3fF1Vmns1nolrcqQ+RA5dSulw6UTEyCkhJCxSm3/6f/u3T//6zb//w/t/47//NDd9pkyZNmjRp0qRNTQb0pEmTJk2a9K70xBNPnJ3TPMKpiBhxNg9nTu8zAPSHCAXNSNU8saWKYIgmJasIgAW3EFAJgQgpJAwRODAFQvZMoNuayACB+r4tXaddxyEQYj5agle6UxWRoiXOZ3FvFucJLJtmVTGOGGYxJDPo+8wxcYgG8PPzb3//pdf+/C+//fW//8F3vv9jNRAFVZ9xDgq1INW2PXPfffc9+OCDjz322NmzZ83gZz/72RtvvHnh7QsiQkSz+UzVKowCwKtX1bnkqoAYEvtCqJjUsWE0EVNzp9r/BLCci68rIiGEEMI6ONUNZf9pzhmgUjJgzbarzgyM57JGLRERCTwiV0oppYx2z7q3papHy861WCzadtl1Xe6z1NTzmtf8y85m/lINaBvK3V3tKFeG3QlS0jtb2XaWd620umk8Flp3usvGXQ+zH/vRTWhV4O3q7uf68vVdX6vZE4A7djvsI2jkZskbJyWK3GjjWx77uzagYTQ6cXjoftEG9ErogeWhGqt6sUHioeqpkzliamKMKcaUkjOCYIBmDO8KrAa0KhJVBMeIf/EjGrgq4xM0QoHMQKSMdCBEQiB1okflO8PwFK9eSuMAHAy457WH0449h949Ziakvm/BzF/EAJV6D2aAVor0fb9cLpeLxeLoaPMc2mhDIwIBMAIqzAPfedv8vnPpgdvnn/zoPR++49b3nZ1h6bV0fdcxYQgxNTMDKGIcEyD7TBg37gFAzIoUIHL6k88iCu5NgxG6E43MFGIsOauqv9txmENTTKUUA2DmIiIiKuK4bVE1MAMKzRwpLpftYdv3pXQF5/uz3B6RLH/zS1NZwkmTJk2aNOldaUJwTJo0adKkSTevp556qiwPLh12t8xDRplxmKWApSPITFaylL63UkSKavFfhYlAVRAhhNA0qYmRQRiRiIGDcbAQTc0ETHXwJEyyaC/t8ih3nZQSY2Ck3PeMGImBKKYYmdLeLMwbniUorZWOCIyCcQLDnEUMSrGu7S5cuvzdZ1/82jeeeeqvvvPqzy4uCzAjICjaug25sjEQQwj7+6fe//73PfbYY48//vj9999/4cLF7z333Esvv7xYLG85e0uIwRN21W93vGn1kcEtY1VFhhBiiGFcAp5fY1ZRU/XMmvM3VDXnXnWNfMrsKT9fTkQx+h4lpeixOObATO7FjHhcREwcVDWXPETSLaYQArt/XUrxlvu+90n0zv1o205KWS6Wh4eHR0eHfd+LCph6QS8A2KjD9Q+v7T7s7NXmwuvDKQBOkE1ew194q6s8OwKsD2fYrm4ZrLMorr6zcZ2aLx3GFq7mqA7I7+tdINvx1eqQrI7J4NpIg4H5WdkBxN1tkR7v4TX8z11x6VWf1qzwwX68elu4sjM3Fu7eyv3Qm0Ve/KKGYY4TSK5KCLrhZo9pt1degc7u2qpPutCcC2LLzE3TzOf7TZOkaVRtNps1TQohDiyO4CQNMzA1I4LVaM1I8XZSh/oQmUvV3EUNIQJAKfWdFkIAQDP05DITaX0jISECgo/PEdH48qzTQNQQYMBxWB2QQ3SKiN9KPv5HBAgQQ/QWDUBVVERNY9TUNMwBAUouUhH5CrB6HuvRIRQDMJBeXj1/2F6B9jDNmls4nZqdOnNmPp9jCcvDgBADcUiGpIZIwb9QBURiZjUTFZGCSCHG0VX3rooKIjGy1QHIEELyo0P0M1LBICLF6zESgCIas98CTjbhEGKICsyayOBASgZZHF1poOtK/Hf/4+984X/99+/+hps0adKkSZP+yeofw29KkyZNmjRp0v8v9dwTTyxONUfzM/v5LSDa2+PIKN2BaQ5gTeBExAAmYiYANpvPYozMJCaAFgJziESEXYdmQGSiIiZqOZdSSl/yGAdWMNECqADANJCR1WIIKSVEghAgRYyEAZEBSobcg2ppl2VxhKGBMIc0P1jkF3/8sz/6j3/+zadf+v6Lr18+XHa5DGhlQAS1la3nciPjtttue+yxx77whd/d3z/VtsvXXz//1ltvXbp4cSy8BQZIGEIQURVLTUIiNVssFqY6n885BFU5uHJoADHGlCIHRsRSpJSc+xyYmMg5pyEEM/VcM5EbItUf8chzKdnM3J7IOZdSYqzhaOYw2nw6dE9VI/GYmfWkc2oiM5lZ13XuO48BQxHpuu7g4ODw8HC56Lq+8zn1ovpua7LdpHblnXf4rVur4c7Vtrc7loDeSq26i3P9poZ11le8oZO22tFGgng9UrrZ/mqlcbRhY02wmjm9dpHDtYTzemfJy8R51BS8LBuY3tQ9MKIurtGLMdMNuyYgDO2s/bVp7O8qtYfIUM+J1vESrCM0Pry1dmV3Y0CO9e0G5SVN3xMZjEbnDW+6tlW9L7aPdmdUe/N+Oz55ANDLFBJzCE2T5vO9wYD2F1F1lnPOqjaUG/S6hcWZF2Z15of/pM4fARvrB66P5cDghgMQgCH6nI9aMXW48Ye889bMhsFxHnLBpYB/pjjySOoQoIeIwYCZmBnQYTBaiiPxjQD8/Xx0tGiXS5V+fNz8nUM+n8EAAciADBLBPOD757NPPHDXP/+1jz98/x133roX8tF+oiZwLyIKYiAKSBzirKgC0qyZwxgPV1NVUxVRkYKIBtZ1vV8fEakjRAZmajXibf4jKaWUXNlKRGEAkgyvCR8LYAMSQCUsuSza7qDXpQILAisE+sKXJg960qRJkyZNuklNBvSkSZMmTZp0M3rpySeXuqSFLG8lDDBPIUXWcijtYWBKgZsYElEAMFUEI0KOTIQGZoPNawZowCImqqpoaGZF1KvwASIFZmYKwUBFCzERM3FEIiAENQ7EISKRARgoMBgBmELO1ne570vXStc3e2c6CxcOu28984O/e/r5v/3W91/5ydtvXVxYhS+gmgGaZyLVbZjBZ7n11lvvvvvuRx999L777r/ttnOHVw4vXrp4cPng6OhouVxyYHcxTM3AauZOIaXkMNO2bc0spYQAotrl7ETUGKNXIJTBlYkhMOFyuUTElBJUS6WgB/YQRETVUkpmmnMezGL0Il0ppVJy13UhRPdQcs6ed3Mfx8+65+ZEpW3bGIP72m5AD9E/6rrO55cvl8uu60pWUfGO3qwH9+51EgP6KuucJLm8w1neOlK86jerJdU+3mrKVtnmnRsDANHIIqi26k6KxbFLgIPfXfECa+yCNZtYEXHLZN/SWPVuFf+1MSw6JGGHPrxHROljJ+vmo8c7NzMzUyR2I1JVwCvgrcEXENe87jEnvqJBbCBNbrJH29Xqbvo5MnkPDGjY5k+Mi7eX6o71dm2KxCGEmBzKkWKMzIxYaxKqvz+gpnKtGqar3Q2n2gxAVEUUsRYC8BXGmRmlFHdQa8gXEQx0KLjqrvR4o+7I5Zu53QyAZoqADuhHRCniO3IA09AaeikCAyulRp7JPy3MsvOVcz+ipQD8KM2z0363oYGPezSgH3rfmYfvv/3xj77/4Xvf/8AH33c6YYDStksDIGI1Q2QOSQCROaaZFZVSnJStIkxsBjlnQFDTvu9XMBMDMKvsdTPDeuOZx7dFzPzjmCKHlNJIsKk3KZABqAExQgxdloO2PywAYBCCCBrzF7/0eye7HyZNmjRp0qRJG5oM6EmTJk2aNOmG9bWvPdEs+Ew/f7s5CErzvTjnIPlQZUkq8/35rEkpMKuRjSEyKppFikg2xIp9yNmKNiFYkdIXDgGRFIwIQ+DYJPYtQ/DMLhEjM4QATIAIIoAAhIaoOZd2AQyABmbW99L1fdcVMQPi5tSblxbfffGVP/jjP/ubbzx78Qp0BcQAABgpEhcVNUVEIDPwlCQi4d587yMf+chnPvOZT33qUzHEv/iLv3r9/OvLxXJvb8/McsljUNMGw8KdcwBAqsjg0TRR1ZCiR5KJyHkXnv5LKcXACHblyhVEms1miGBma1PIq4fjGOiccwgBEUSUucJY+75bLpchBOeytm1bSkGEppmlGEufHfyZUlLRxXLhDrb3zZOALg8+Hx0djVFCX34sh/jL1ba5vO3zvqcG9I6tbO1nxwgIay2sBZK3+rJmQNvxHxFXNIrphm12EpIy4ggWqFFfxx34zohO+i/esQUAWIUj15bbCCPGXWf72rKdWPUToaJPqFVaeXgqPdPqlpyKmhkx+XIA8Np0pnqsYzuHWm7agMatDW9+LOcfqQFtlT2BNJb7SymNKCGoLGMcRhXrbAw18xC0B6Ldm0amIlpKORaC9qa8iKvvYTSIPa0MzpVG8FkgZipy/Dx7grgO6qFXPURm5sAI2OdsNSPMTISIXs01xggEDoB2kIWaIQBD5YF0ue+7LnedSG/18wMAgcb4uIEhGSKZJrMZwMfv3v/0Q3f9i8984tx+TJZzd8RoTQpYN2bjgByQQu763HYqoqJgFlMDgDlnIDOwXIo/6TFGQgQ1Yh4ZI8OFt5rENyUwRGSiGCMY+GeMjwn755+ZEquCLRWxmbUFDjtQBZtF7bMV/W//tz88wS0xadKkSZMmTdrQZEBPmjRp0qRJN6annnoiEHAEvCLENm8Cg0G/ZFRGRbRmNuPAoIqiaNVNZua+70QLIvCA4FRRUJvHyMTkFlEI1jSoBcEohjornhnATAWH36gBAEChZDA1U1HpuuXR4SExMYcQYs5ZRGfzUxhmbYGnn33ha994/s+++txPz7954fKVvkBRUANCZCJCLlrMjIkMzX8dJ+Yzp8/8+q//+iOPPHL33Xe/+OKLL7/88iuvvBZCmM1mJZdcsoh4ahhG+gEgcyBiZyUrQIwRAfqczczAvKSV1RgmDGhUMzNCcJ8whBhjXC6X7lOPEVfCVRjQU88AVkSYRjenEjcQKcboLTsnOnAw1VJKyWUo2IWqtTikRwsXi4VHoV2DJe05wX+o4HMVwvFagmvG+FiO74QG9E7nenuXx1fbzCPjepW69UZGgu1gJB1vxLfYlbj2TXGwkuGYE30NuQFdWxkHRKyWjyPCMeJ4nXZow4D2PqgZV26vW7XmXvnNGNC7uNDbx3Ij8WrbihcDjEaqgZk56wYGA5qZ1dQNaCIiJtPjNuVYD29rTzcl3eCHv5uMt5luOMLX7dJO/rXVwYSrnrcNnTABPe4RvPYdEYfAMca9vf2madyoZeIYY845l4Lja3PNgMZairOmof0NGUJAJICK11cVLxioaiFwSml8UgZnH489lauDUTXVEINDnLx2a0wxxkhIOWdRMTMGrCyOIog4mzUKA4ZmGG1EAAZC9Dp/VEpul4u33nqj61of2DMzXE/V+41tFgySwZkZ33Hr7IG7zvwnD933yP0fvG0vsHbWL+ZNIoJSiiILkBnkPktfmNDxU2qQRfuSAYECxxhDCEzkz2mgICIqauBB//GpM8Ix3g9ogIgmIiIlF3e3Y6zcrCKdWAGO1uyp8bJoJyBIKsZM3NDvfunf3dhdMWnSpEmTJv2T11SEcNKkSZMmTboBfffLX17osoWeWwgBm8SJRPqlSptSCkwVEeu5WSYCYCIgZ1wgERMDIRA4EoAJIHLwunkAAEQQyIQM1P03UJOSzdTMQbqKpugsVymIho6HLjmQp0fVFDjNiCLG+c/PX3zuhVf+5hvPfeM7Lz7z/Gu96DBHusrMFNxYQDM0MGY+deb0hz/84QceeOCjH/3o3t7eT3/605dffvnVV19bLpdnTp8JIfR971UEfdbziLkYQ6zMTEwG4PzQhqjOkqaaO8RB7lOICIKip9iIoFbEshBCNTIQa8kpEf+6xpnNKqV3iLtKkdHgHpODzAQGRIMFgUBEquLUjq7rcs6Hh4dd141zzMdGbpqG8K51LRcSb7pbK3vr2qvthGyswuC2ZoCvnStYWX03Guyt2I2VdWZrGeTrb6115xtOo5nTCU7onm6nYqvTBzJ+CwAqcsJejQ2v92e9+WN/w2hAn/jk7fTWbfUz0AJjAhrMxBTWD6S6mWNUdbtHUG+3d4Hg2NryZKMgu3VszWv3amM4YbXsPX+m1zqlZqjVKVa1EKLTfWJMIUQOARE5hHo+h7Cuc4rMN6/kjWpAE7EPoljlbHgZRBgRHAir/+rr1BPOdHzgykEWHAIhmlnOWVWRsElNCCHEKCJmGpDcRk9mhBRjFFUxrZwcc5wLMBEYOCqEmRBh/9RpJCy5d8DIcB/64wzu/QtAb3Cple6to8PDRa+h7eHR++5436kwj3tFivV9yb0RARIhQSkq2QpCCBRTyUVMkEBMQRRjgMqHNjEFs5JFVIcdm9Yeok/KAUBVdS65DVwlAwREp0gzEzEjIBKrFiXcTwnasiwQiKlBKPb7/+oLv/u/TB70pEmTJk2adAOaEtCTJk2aNGnSSfWt//AfoMFocZEWxNBACdaSZdCeQOfNPIRIRGqKhDHFxCEyB8QiJedMaIRAjCaCpggYCIdkZc1wgqnl7JXCdCiX13VtkVLnNQMQGII5oCIECpEBjJljTH3WomAU0tlbeH7q8J3lk3/y5//nv3nihR+9c+FyawxZoazl+apLuxaeNbT9/b3777//t37rtz7/+d949tlnv/3tb3/zm99k5sCBQ9zb23O6hXu1zAwGOWdiCiE0TaNiqjafz0OMxDQk7JKbMX5+VLRWFiSf541mZipgylwJGyNYwx1hM3NKadf1nsJeLBalFB5gpqusNIBXnBrdDy8uSIA559znEAJUorT0fXf58uWLFy++8847Iw9kQKmOzI1/kH8vbcSZd/iRuEbEuKEE9AnZEVsl+9ZJEdvUiHGJnszbww3LdTPcPdpWuxzP6zrJO7DFduIQ61acGIkB0VTcLkRiADQtV9l+d482vPjBdlxZujvT2SfGhlxLDpznWoQQVN22BKJ6fc1AZA2fsjMvP4aIbzALXLfadXRIx8YnTog0sW0Ex84E+NDqtTpvQ5m6jc7eVAJ6R2jdQNXJMv5inM3mp06dbpoZIjZN4282G17yhBhjdI5zUfUI9eqZUvWBNB/scX/ZCwL0fX+0OBr59V75sO96IoopbvfUX6c+XEgDDKrv+/l8nlISdbqGpRARQFTquxMgS/Fvzbz8YG9qwQsnqnfJAKxIOTq8cnD5kiP4N0/RGOwGUGCAANAgnI7w4fed+o3PPvbJB+6+9/azB2+f7xaXQfoQMMYwm81yLl3Xd10mjk0z70tvBM286fpORJq0Z4Aq6rhtUbHNoqf+2RECjfN1pBRT8/FIQWnH2gAAIABJREFUAh8PRkDolh0CNE2TmsiBRbMZKGBbrNfQZluqUSAz7OPpI9r/qX3gS1/60vVvj0mTJk2aNGnSZEBPmjRp0qRJJ9RTTz2RSmzakM/qPPHZ03vRiuUFo4IWMG1S9DiYgSECE4AKqqKpSFGRJiWPnWnJKuoMDjB15AAhqqjkknMWVTGzStwwJ12kZkaBAaCUElOKKVGMaqolEwM3Tdw/JQXNGLg5OGxfe+38k0/+2d/+3Xefef5Hlw/7thdDUABZt1hGh2NY9OBDDz3++GOPPPKImr719tuvvfbapUuXuraNMTlbw+c71+iYaozRzLqujTGFEGDwmvxXffRMGdgYahaVIZdXw6qDAweESIQhBJFaV8o9FzMjwhij0zlF6nL3ix214Xv0QyileKW10US2Ic7sEpHFYnHp0qVaZ3DpxQZb1VojbNPifG//sbQjVrwjz1lDyjt2vWYQ7sJYAK1b57v3g7vgtzv6tV2yb0g271pzdd62zTifBK+DkUcDLGM8xqtEWh0r7nBWh37ArlqCuPN4t1rcAb/wAYbaeTURn5lwfCVEMx3i2QAA1VtErKgBBc/+q0NjBu/YDGrwH9Yr/flVrI6r92x11QjBmTReSo7Q8bTrUfxrBuNXadhhqAFF1QCIqVLVfa7AwDlBxzLY0PbxCzKcj/VM9XBlhhEaG1bbuid33qS7yRknCn1v46TNp4PUFq7exLZP7Wf1WCB9O0q+9bjsHgLZ3nM9LUiERMzMnjIGwKZJzWyWYlQzUZEifrm9cVXzQLFuXpSNvSEiMnhxgFL8ZTsMtIGI+qDcVserxvez1ZvN2RigKkzsLrY3vnHI/iAAImLJGQCcyD/AjnyoD0rpu+Xy8sHldtmu5grQEDtH8CFUNCAABmsIzs7Cfe+/5dH73v+Jj91x7x233roXorVWFoxl1iSkaMiqgMTE0VANwdBURUTBUIpKlnq6DGNKgQMSShFVQSTnyvsnVxEZOlLxITzUue37rKZOxCZCP2Oi1vWlYCxGnWgvAETM9rfyyL1nfrL3oYMvfnEqSzhp0qRJkyZdXxOCY9KkSZMmTbq+vv7kkzn3feztFEfGZt4EMpTCjAgEGBCAmE015xwDI4Jk0dKBFEKrZi2DGJqKSjHPAksxFfBf6M20iBYptS4VAlaTiAPH1DR7c4rRAFEkppRSwphESsmZI9NsBnunsHC3lAuXj154/pVvfuO7f/gnX/3hKz8/XIi6j2JmOCQvh0NzFzDEePrMmTvvuOOTn/zEgw8+eOutt770w5efefbZKwcHiLi/f6qZNYGDiIXAIQR3kM0gpahqSJhSYuZSiqMwEBGdM6L+W7wikkN0EZmpRtX6Po/OiQclcy7OZTZP1lnlODuLo07r9gngYIiDwbcWFRQRAAvEWC0GLGYi4jk+A1ssFpcvX75w4cLR4VHbLitzw9woWTe43vNx+qtlPDejoCvHa9fKGxbbMSPMTcdtYjUObW0Zblfpw1U1DheMfQVYQZdHP3er7eq/jkblmPpfbYArVxLX/kbEkcGNCIjHosE47nVcstOFRCdM19vfLVpCqpQP9DkJCEjH/WdAA0DbNNmJsHq9BgbAQMzu4xHTegdQ1HdnZqMxPPQT/HD8TvdFxARq/h8SEZOKwlBibh0JMzyD1UsjRFUzMBqKMY7dIEEA2KjxCDY64AAIoyu9ftibJ8LATG1s1O3ctW/8gm7deDiGqjfu27G46I3rOBYHAQ1pdReNizfWgu0bs958G/3CXc/Uyfp5tVEdMxVT0ZJzyZkQDSDF1DTNfD4nZsP1UqumqlLUA8rrBIsdDxVs+MuIQJ4r33VmB+dZRyrRYDEbAnAI/hoEsxBCCME2NjJ/CSOhytA3VQCfR6JqzhNHZiJGAAgphhRDkVLH/9ax3X4kaIhioGCqVhZ5+epbi2V7tFz2Ag/cfe6Dt55N2EToGDXEhuMMkBAJvBugWTIigoEWlWJa6klEoFQNaMo5uzsPZmrGTKqWcyZCf9V71UgPgwNBKSJDBcURxW5qzH0WVbPT+/tdtsOuF7TPwPcOPgThe/DEv/yXX/y9yYOeNGnSpEmTrqMpAT1p0qRJkyZdR19/8kklI8UcC0Wb76VEot1hMCETkRyII4cYqO/bo6PDM6dPxcCl76xkBJ01kRBNlQhNSu47MGXClBIOc/BVteQMZkycUgopcozEBBwgMDBjiBgicARmQ0ADVAUpAGDE0DQYE3DKHf30p2/+1Ve/+cdP/sVX//rvjxbLPmux0SWqaT6FtbAqACKeOXPLY49/4nd+53f25rN3Ll38+te//s7ly0DYNA0AlFz29veIeLloU0pN0+gwU9sDyG3buqPhs7lLycycUooxtW0rIh6p8/wykU+Fxq7rrlw5nM2apmliTB7la9sWAEIIKSXHNOdczCyl5Pafao3UeeS573NKKcaIiN5CKcVUyeOjiIhYZ50TLpfLd9555+DyweHRYdu2IkVVt7i8V7OJ36Wu2uym04cAeA3mx5a7qmvLt+OhO8gGhlteGe6Ijm7buNu+lg8dqEjlwxAj0XaIdAUghpVFO6aPYXCud8RiDZCQiUQrtgXweO99CMhxuzBU1TvezpixhxV8HGu02UTUg/m8RR2B0YTzfY1/Dkl5VSGiwKxW11RVAHNSAQyetQfwCdEtMB2cPUBgZjVzZC0NkX83/XwTNTNRLUJcYQi+ixijgYnUDUPgnEsRWTeg/bQ4kH19TsB4NdcO7jpSVcmZKh7XazOuTtGuLbBeG4StIG4th3iS/R7bBa1M72OUhY1HGLfX2kJw4I5M9E5ayPENb9Y6H58pI2Lm0KQ035vP9/diTD6c0Pdd3+ec6zAeM4OZ1KkZ9Y3nd6y3d6z57T3S8JSNXPsR7lEnlKgSUorRV6i7GMx6q7hwMzUcWEnkpQyGIxoi1EAEiCYqjkkxNVEpRXLXScnD6R1Hm3B4JSKCMUgCmzOdafjjH9z/tcfv//x//qkP3TY7ncry4CIzh5gAEJmISURFS9ESYgwc0JgxMAVPLKs7/mYIUEopIggQQoghGIColuzOtT90wzAv1tkjPtBSXXcwR0X1fS6liAryzLhpu3LxytGyLwBw8D04+uDpV2+5Z2JxTJo0adKkSdfWlICeNGnSpEmTrqWvfe0JWfbcpX6mGIxjtNJ3uWXLgmpQ2Q7EVKQA4nw+5xCIkUKkEALjrGlwmCeOZs3ePpgSETcNYqWympmAIRgRcQzkhhEMeU+fHS0ZwMAIwUDFpGjJaqBAZRHbAofL8q3v/ODp77z4zHM/+sELr1x85woAKqwXoRpBBIbVg9AzZ8/eddddjz/+yfvv/wiAvfaTn7z+858vlm0IITUNEbl7m3MObF4DcLFYmKmIlCIhsKr1fT+YGlZKESkA2LYdMzsDOqXkYTRwLyBGROi67ujoUFVEJITs6Gdfh5mXywURhVAZ0EdHh4OnVjPjzAHA+r4PIbpvMlT9Us81+jRzJm7bdrlc5pKXy+XR0VHXtrmUYeL4NtXgpt3nk2y4vc4xu9ntGbSrwAS28tmDubeeKd5Yf5fxveVcbQVevbHrH5GZEdPYDTMbk4Nr7dAqtoowwm3NqmvryJQd+yNEADUjJAo0RCeP9+AYg8XhLdsHM1quNU1MiB6NVNUiiAi8w1j09ZEJnL3r1HIAD+MDOEXZw8cACIO7XEubEZO70oioAJJ1YDrUHmoRQNBqa5vmDEiGAGpAqN5tNQBQUXUzdLS/zdx2B6ZrRIq9rBwxaylmRo4SHgg4ZtVbXB3v8VNQlyOuvUwQd3i19SdrQwsGYDByHMb2dqGWryUcw/LHF9UWN7/bWslgJLfY9jO0Y8P1Zdd/Dk5oSQ+rmTOW3CntS2maxkfROIQ5h5TM34TVF2U+ZkATSR04u56GcRZy3ohzoz1b7VwiIkZEfyoBQU2ZmGl8EobXi+06CwgIyH65cd3NJwSjgAwxJZDUlNwvF8th7HC7mqUpoBK1arLMPzh/2NNPDjv5Z7/y4MMf/sBec6tBERPQEpA4REQDBANkQDIsfa8gSgJ1BkwR8QkESPVxRUZAMCl1xJEQwAlXZk6tV1zrlZlzbwwMCAiQ0Yz80z6DYArxzLyRIp3q/OP2fLjns9/72o6ZH5MmTZo0adKkNU0G9KRJkyZNmnRVffnL/zp3Gud9B8AhpKZByaVdsuYQkYkIiUJIMUQOUgwDx7iHBAjGxBw4Bm5iAjD/vZcJY2RQBUKIEQBAxUoBBAxsaLAy70zVwBRUTRVKsdxD5cwWNDXnRYtlgUWnb108eu38pT/447/42289/8abi76o1ejhZvpwgAEQY0zp7Jkz99xzz0MPPfT445+YzeYvv/zyK6+8+vbbb6cUYwyI2Pd933dt2xUpIUQmLkVEylCHKhMRgJVSKoC0xkJ1bZa9p0G163r3qWOM7ojlnEuRvs9mQJSH/KiagQeZiahpGqdq5NzXCdbVEsK1XXdEqOp+glMCEAdGgYoeHR0dHh0ul62ns+uYQY27brjz70Inz03v8KCPf7uDv3y1lgbfEGCdujDKKnjiuMl9PGS9BbrdbupqPhwOhrLf5DvC1FTDxjVxPwaNR56wT4av0JT1rqM/OzQSCbZsHgMAj2dS7YOKupt2/FS4I2o1gYyIDlU3rRa2mmI9PetbGQAw1uQp+SM6ZHjdXxZTVUPAgf7s1IHqNrrZVx13FUAEIqyX2Bw8DbUnakWQ2UnQYOh11XBwnG3k23i62cwzqqogso1eAeeEqBQxRK+uKTLa3yOWeu2UD7bmZrq4toYVh2JrK1zVBl3BolcW9rjJScY2dghX+z02xLG18zVEB2w8KSsY9A5DddcUAoDrvhxwB/fmWjLzWLsWKW3XNU2azWaz2ayZzVJMIbIz7r1lQhSz6hEDQLVZVfVEeySiwKFnVtUYgmfhRSrdaABPaw1EizBzDHHAT4/x4JVU64wBP4OOrzDPxJsysbfMgZ1JbWY596qQ+161mGgdlxhPhp9AJAETtZ9fkYMfv33+jbcNG7V43x2nTkWKkLVvmS31wT8ncpEQEgJ1bedPCgCoz7IRMQAkbNKsSQmJpBQz67pOrX40I6KKqNYxGAUzUBzo9D44o2BcuHAQKSKiIgpZoVdjpnQqhe6oA7RPwzP/5e/96c8evsue//nkQU+aNGnSpElX0/QpOWnSpEmTJu3Wl7/8rwNQAd1P+5F5tj9vYmAVLB1ZIdLIGAM3MQIYqDEhoQFYkWyqiEjovEqPWmkIkQJjYCgZVIHARKwUEwEEZCruOYGBmqmCiud5VVVKkZKRUKW0y0UIAZnavnRZl538/I13vvfCq9/49vPPv/zmT9640vZuMmGgBIbiIS8wAwEAT3xR4NvOnfvt3/7tBx988OzZs08//e0fvvzDCxcuuKmlqlynHvc551IyEftv+M7PMDMRERltCK+axTFGEVWV2WxuZn3uCYmZmIOqqHoZKFBVBwWMxQlzzk2TYoxt2+WcRaVpGiZyqwURU4o5l5xzCLUnY+7VhtApIhJxCMzEgbjt2oODgzfOv9G2bSlFVN3g9uuLSFsz99+NTmhA78wj35QBvWpph++MKxTsjj2O7vNaQNQ2l1wVwbGxvCLF10x8BNsKU7vjbDKUguTNBDSAl92DzQy0jXjeNdvRDbnjB1upFuuLYMBTD6bnaD8CwGCAIuKABEBTMRHnCGw0XisBqt+u6iUBDTxfaUOMcmR6kM8DkOINq0h1YlWRkJnH9of6b37gI6BZibnukajWT1MDtRGmssJQD197fFxlBwPazLwQHHlCfEyAD13eOEtmI9F7PQ+6Ondr5+bahvIJ4/PXXed4s7uqGm7eNrti7MeOsUKVt2g064c9Nj40cJ1dnOhYxjz1xrgXEhExh+Bg6L29U47UtwFwb7Vw6Hr3dvB2YOtUiCgTpSaVUsAgNY1X7pM6j4SYCbxwK9RJCDW+D/VhpwFlJEVU1UsdjLAOUWWnu6AvFgSQIqXklBIxm9YdlpyPFoeLw6Pcdyrqb731S0ljDt8gos5IPnjm9AMfPPefPv6hB+99/523zY8uvZG7Kya9lxAoRdC508jVCmdmImb2zxoDnM/mTWoAQYr0ue+6DgCapokxErH6MJGqqKmpggxg9OHBQKxB6XruzeqQHhk3imnRlV4BAmqk/+ZLf/DiP3/o43/x/RPcBpMmTZo0adI/RU0G9KRJkyZNmrRDTz31hBXJms9gExpoZk1gYhVGYDBCJVBEI8QUqp3Gdd655twBQFMRz+qFyhCAQ0BPWZrW2nxSVGSwAK2YGAABlD6XXMyUQyDmXLKq1ZSZSs59SIliU4zfunjl1Z+88fVvfe+73/vh8y//7NJBPmpF6uc7MQao1c/8l2gxMGKe7+3dedcH77v/vkcffWx/f//w6PC5Z587f/48DNgKqEaGtW3rXoOqIaKTms1sNpsRktZ6TW7MKQA0TXL/umlmBlZpmyt3ZrTpfCI5pZT6Pnuk2sHQpThQ2OdOExHlnFU1hGCmquaQXHFPjZCIYUAJ+LTqIiX3fdd1R0dHBwcHly5eLKWMYdTxEt9oaHFT100x71yyayFusy/weG4ddmQ8143lrTJv64Xajic4t9xngAEOvkqK7thbrSNIg//r55sIHSdQa+K5f4nVzaoQhlrLa7D+iQbmc3XfzIvgbZJABqd0cFgBwWERRKZjiHUtDKy2HmCsidHhwLWGGqtV7Igb1VohEAgd4OKlM8eTUPPciKaGCIikKmDAoysn4isNXJFapk/qFP5199ZZPbzuhJoZ1nKGqDYURKT6hMDwqIAB6LFyeU622HAzx4T46giG0+PLmRkBRvOxjgcgOhGiXlMwAIhMZ2bxwmE/FI+0lXG93otrPkE7PeghDg+37cdzp5t55CZyZMxifZFFLxeudBcOO9kV78XhTxzMd6sx+eP9Wvv/2glby2T7WMn47h2PZxdXxI49QttHPZ6768ldXdi4ZMM1Q0Rn38/m+w7l4IGXr0NMeP1kOO1mfdjGSS/1zWYAAKJKiCEGKaKmzGFE1vjDtnpkBsf52AHWnhGqqJh6onl83tV0/EJN3Z1V0TXuv4+qKID2fd93Xd91fdd2bTe6/7i2I/+CzAhkBvC+U83H7j738XvPPXD3rR/6wJlTCVg71GyqImoKCBhD8s/eMEiklCKlaIwxhmiVs6MyjFkODjN60Uf1op9g/jYgHjHZgxu/dRVVUSmqUa/aCiECRv7QN3/UHCwf/OsXpl+wJ02aNGnSpG1Nn4+TJk2aNGnScX31q/+v5KIgnG0v6SxF0g6kRzMACkyBkQlz7lUKojUxpRC0FANFtJJ7Jjp1ag9MQQUBCMHdKS0iuSNGQkRQVTHQwMEARKSIAAATt4tl3/UKNN/fa/bmbZ+RMKUoqoaGhJT+P/bePNiy6zrvW8Pe59z7XncDjUYDaIAYiLFBcAAgzhIlirIoepDssijJkZOKrLikTFZJLqdcKSspuFyuVBL/43KqEsVJpWKXrCpqiESoKEKmBEkEAUIEJ5BoYiAxNIBGN9jo7jfc4Zy911r5Y+1z7n0DGt1okICA85EFvHffueeee6aL+61v/dYYwihb9ejjz97/lw//f3d/7puPP7s+96gomgciC86ji3SBAQogrqyuHjp01R133HH48OHjJ04cfe7Zo0ePmlpd1/v373d/ucspy2w2Q8TxeMVpG3tW906n06ZtD1xySVVVAGCgRMgcfNhgXZdRgUQMUJwOEWmaAolWFWdAp5Tc0Z7PZyISY+XwaCKOMVZVnM8bABiPx03TNE3jHnSMAQBylpTaGCMRiSh3nouIpDatra+dOXPm1KlTm5ub8/nc7ezX+hzZJVa8wwh7WY7zjjXtSEDvdNWW8buLJ+5Ia+54xdU6MtHmPPWO3s5lVmq+Yv9oFPnI82vb/tSnnt0Jxd4+NnACADFKVgDg4GlHR1EgFnb5wnfepusuXR1HOr4232hNVBb28fKrq5lZJNyzUk1aSVlL1FfLCLwyz9AK8oIDg7OSTRHQG+2Z8M5r96/P2o15mjY5q7VqCqQGOedtZmLxzbsdbF0oGH1om49xQ/QLhBEItGaqqzCqY2SsGCNTHbiKHAgj4TePrZ/cbN2ws07+Qu97+yXjio+tzU9N0vo8JdkCMMGlsLY7tv2m+hEUyQA9X3vhG26rshR0CYCZBWZE9PtMMabLD8WARoBL9tTvufrif/jRG3/z/mf+6Bsv+OPiwOCXt1iXX3RXV7qO/N63H7j92otvvuKiGy7fc+memncc7qU1wJlp+9yp6TMnJ48fX//60TOPHV/3883ACNHnTHbslN3Xs20zth/o7X8sJaplH7lb5jUaQli85ld4LiJRCDHGGKvRaORsaFEBRHdOfQNUAfrcfTce0LFFiM4jAgRw85QQvWHF/WgH2vhuU1E3vtW0X5iJ/fzb8k4RDXfZq/1LFwt5Z0Tdyr3Qty2nPN3cWDtzyrq2Bdx+Py3lJgYIABHgygPVbddf+lOf+OHD115+cY3WbGpuVcw/D0NgL7DGGAIHDuxkp2be9HY8EYUQPLXtfCdV5RDcmNaSbDYV9ToNE4EXtlQLWQj60g6YaLc3Salq2jxpVchU7G//yz/43Cf/2hfe+UPDTMJBgwYNGjRomwYG9KBBgwYNGrRF9933BybGMdgcAiuAaWpAG9AMAISMgQBJuxCmGaQsYIZoKjmn1kxj4Da1oGqawb++moEZIUTCnBRM/Ts5M1GM/lePjCFg5KB70GLkGDiGWNUQmJBMMqgBkmJ18sz0vge+9Of3P3z/Xx45duLkPLu3Ub7IL/XMe7pNPMX49muvu+Xw4ffcfkdK6aknn3rp9KnUpisPXSkiRDQejx36Yd3IqRACEdd13baNKhDzaDwOMZpZ07amSowAlvMUABxQIJJSSkSsKm3bumNJRKrikWdVnUymZt6avVFVNTM3TeNbqyo5o1tCInL69GlbQjbnLG3bmEEIQVVzlpQSqIGZiGxsbqytra2vr81ms7ZNOScAw3742GtG2zgX7eJQn9+ztz3QoyGWg51LOeKX0y/96I0//+HrACCLtVnETBVETc2IMBCOK45MADBt5ZP/5i++u9H4E62brll+6Z0+K2lJ/5dkIyYEkJSQkJiB0HmyoGVRpO0xb0L8X37ujusuXQUANWuSNtk95GKBEWJgDIRVKHnpX/i/vvitY+slNYyIoViQbtEyE3DZMxyYgXuSwJ4q/uu/f+fOPWMAopZFszodBKyzxLBD3zKVWCYhEpWwMvVZzXPQr/zmV09NkpghAgLmbkCiin7s8GU/dedV/ZJJtM1lY/rQ5db9tsAvbP31FbTzaV1gvo+9GxMGppWKu3mRICo+ERS6k053CwifZU8gYhXoY++44m+858o7r7ukCudGNgdAhP2r1f7V6l1XXwxwFQBMW/nK06fue+zFP3/sxVOT1mse7mmavazXfJZLw3Bn+WaXZWCXKs+rFb7s2MYtL2qmkhNAfxOGLjauak6rEdGOBwHQGcX9pVGuNnMEhxgAl+6EEpGm3sU2FVEAcNhRufoICcnT0WXJfrDnTvpN5/CmnLHwpnnbxe4bysSC2a9KjvVFF106mWyktsHu0xGXnwEIgAKoABn0+EaWZ9bq+742nd36kfe+s451pa2mNjJFIjALTEyk4kl/rGtcWeknE3R3yVL3ISLKOakKAPocB+/IUbOcs4qUtL8BYnGrHUhF5IMIVXJ25xoQjSrhuDpt1zZnc8h/+Ot/68vhvR/55n12QR8AgwYNGjRo0JtQgwE9aNCgQYMGLXT//Z+SnJGDNBIqHoVK5ptimZgMGRGRGDlSIABgJOJgAIQAhMzEKkiMaEyExEiGEMBK9z+YMmGIrCKgAmjoDdZVBDPwuCahEQUgIIYQ/Cssj2ojNFOjKBmaZM88d/zhbz312T958KGvPf7Yt49t+76//K8O6wl79uy57LKD73rnu2688caVlZVjx46dOHFi1syJaTQaMzOAtW3bjwH0zGvOQqQA4JGxlLJ7IpPpFADAjAOpatu2zGVwlift/Cn940RoBs7TyFl8GqE71CsrK8zBJ265WUDkDiSmlKbTaYzRiagA4Cs3t/MQVS2llNuU2rZN7ebm5sbGxnQ6yTkvvJsdTeWvkZZXiOfw885nnUU7ws67kQHOreu/KDAGPtt/+K1U/Ks/cfif/c7Xy2tum77WG3a29QxbbM6yidSN4HMOxo7d8Mn3Xe3uMwAQ4rjiccWv+BaIyImtC4p0gVYU9aYSAJhatnyWtSFAIAz0yq97IXpxfe6AaodHd9ZW99OSIpNXAt4gMjUTXWqlKJHbhYMNS+fpjjNx37j6T3/wuk++75q943jhG7NS8Q/dfPCHbj743/3Ndzz4nZOf/spz937rhBkQo+mWHXku7vNi463b9v5s32747zJUs//by/12YTJTUJBsAGYqkiVzYUtE/3NXGMACeSmVG0MkVZX+igAQ54KbUdcMA0uxZY/xGhgY9wa0GXZZd1nwyp0Vo1t2RYlfE6qBSllYd1RnCgGGUU3VI9jIoWYRQcCcWjPpk+HdYbCeCiQAG0nlzOyrjz7HHENVv+3SPQdWwwjzSkVEkNs2EwZmn5hgpiFURARm6jM6vXKMwUP8BmgqYIqEYIRGbrczAjEKgPi8ADACYlQgZUIiIyr7mwKAERgBgCEoweiivRzo1Om1bOFD+csf+53PfeOT77n3nft/9K4/ew3PjEGDBg0aNOivtAYDetCgQYMGDSq6997/p21yVUOaAcdQ15VaphiZApKBCBESM0YmZiYGMHAIMgAjxMiBkLBzbiTHwDF6orBHYoCTOMp0KUJAgNx6ONpyNkSsqzIJzRSygAg0jWnO0irW04Qvrbd/+B/vu/uezz/y+ImNzbnCsv1RXL+Fs+KDz4yvuPzQj3z0R2677TZm/tznPufJYo4h53ypzkeBAAAgAElEQVT69Om6rs1sNpt60o05AICZW9Lm4S9Vm8/nMVZVVfn4Qe9UVtWcs7eHt23rnc4pJZGsqlVV++O+ff20uBgiAIhkR214B7dDn/2NMHNKeTqdrqyMR6MRETdNk1Iaj8cptRsbGyFEH4e4ubE52diczqbuTff2SmlNR+pciNdQ2wwnXPphOcm3M8m887m7afuALigt97DE4kDr4AAd9LdLI8Krtd1//LZDv/OlZ7/6zCnwk7ObX1eizWrLXfm9zaSiAIAczMzEweBdgJqYA6vqMohjTx3+ix++4bw2DHzCWGCQ8nJnV4esMPLc8uunF05PclZTExB/RNXb/On7Gch/FSqXEkDfQ0DFqStYH+jCreD3PCvPYqKf//B1v/jDN+wZvfZfNJjwwzcd/PBNB184M/vN+5++++vPz1s5lyfuTGqbLY+57P69I+FtOxAcu+s1K3E5A7kU29q2pfk8VFU9qldX0OtwqoJIgUNnGRuaB5m5I21I4FAgRSqlCwHJC4EA4HP8kBAgAUCM0XE3AGW6pld6Olw4BmYg3ObFY8+HNjNmX9IUtlVWtLjkZaBuCAHJDGG8ssohrJ05U8qzjuxZELetI18AIjRqz353svHgI996/PGPvPfwO6+/7KqLqn0V1JDmm5umwoQxRDNrc1oZj6tYAVjKOWfRDOPx6uqefaCcksybOREwc6ii11uRKASOMRr4yN+k6oa+n+kmguqgGypdCYSESACkJiQWYty/ZwzNbH3WJNE//vWfrMKGCN9710cHD3rQoEGDBg1yDQb0oEGDBg0aBABw9913p3YSq9lsPdQjHdVUBWTAUI8jUyA0yR0Dt/TjMxFRICQiIAQEYwQmbNtGVYkZEU1Nwcq0JfMcpHQOon/BNixRLWNnFaiBChAAswFozrN5m9WMeW1z45EnnvvM5x58+MiTTz1zsmmzewBEBFC8wm0BXGJaWVm58447b7r55iuvvOrII0eOHj367HPPqmiIARCIQ4zRIcsiAuCzAVFEPPXsTiIAqFrbJlUTEVUlohDYeZg5ZSJvdi5gWR9dOB6PRTTnrCocgvsjhfWMSMRO0jCzGIPDD+q6djy2t0t3AWpyQshoNEopiSgR5Zzn89y27Wwymc9nOUvXgU5OU/B94Pv2e0OCXtYOkOlrtdZiN9Mi1I69jY2w+Gf3jHOFQ+z2agj/5K8f/s9+4wG1EmHGUg8AVSVHiVsxl92I2Wm7FS+cCQ3ALCdPay6W+4c/csPFK+edilXVnLIBEJOZhybdqCcAUBEr790kC2DhRzsT4NXsi9dCSXSehIm44pTEzPx8BgBAoAs4Ut8HYSEFl+wzIBgY2nJ1q/9n2fNm8PaDe/75T7/78KF93+vNO3Tx+J/8jVv/8x96+//xp0/84dee78/Dcz//d7Okd72Cty+3td63pR5zQZ0Wu225malIauYmOedcxRhjZGavrlG5Gfg1B4Q0XhkTUtM0SBRDUC/+dMMJmZxTYz6TkJhGo1HZ8gLUBq/ZOL5my3tG3FZQ8ye6qZ1zKremUpPd/ja8LQYAiBnBTDVWsR6N6tF4Mp3MplNJyUz63dq9BgCAGiS1bKAza6W9/yvPfvf4mVuvXXnPzddcc9l+QIbcgGYwQ7U6MqhoThyYwAgMCVRSM53mrCKqIkpkgbHr6dAMbYa2mfafGv3RJCZCaNpGclYzDgEJVZWIkRgAVUHVANcEuMmCJiCQVEXG43p2TC6/6667Bh70oEGDBg0aBIMBPWjQoEGDBgHAvfd+qm3mTbvKYHWVx/UYdQ55TsyRKh8spsTQDyMCBVEAIqJQws0mkr1fW9JcVZBZFM3dZ59jZk7w1K6PXUVETSmyQzYrYiAGNdGUTYXQUpY2zRuZCzVKR544+vkvfu3Tf/QXp9fnrXjrMDqs08y8Y9oHv3mzfFVVBw4cuPptV99+x+2XX3b5dDp75ugzTzz+BCLGGB0GwIgxxqZtzYxDIERmrqpaRHo32XO1ZkZUvGDHfXJgVSGjkqdDZGZ32Zk5xjgej9u2zTmz56KZTS3nnCVxJ/ediVBFDcBTe32QmZlzzqbKgRFQVdtmLjmpajNv5vP5vJm3TZNTKlm1zi532Y6xbK+RdjW5Xp2fuPNZO/gbnrorVtMitGlAizzy7i9/3pt08xX7fvq9V//2l45CF6kuMVczIChxWCsmc3mNBeykwzR0sUgzA7U+MIsAV+1f+eR7rz7frQJPoqoiIRGbOtbGkJgQwfkWahQIDNTULSwiIkbC141rMWnEdwsxoygYdPAQM305tsMbRT7rr6PhLjxoMFxk+5ej/4AfPXzZ//h33rlaf/++XxzcN/of/s67brnyon/1mSPLj+PS+dm7xK94H3Ba0Za1LF1xW7SgZ/c/lM4D254A3rZdZ/1L2bVbnu/lllYl5Zyrqq6quq6ZgxGFyABopr0XHWMMIfh7ZaYylrME1ZGQOhJ1i4YAGEMkQhHtd4/vtkKLdpqNmfOOoWuwgP7mUAxoI+82AerJ1P378tKEY0O8pGGqXpIMIdSjERArYDubSk4qGUoUerG3FMA7KDRDm609emp9bWNjurK678Deiy/dN76ogkTS5tSgaSDK4k56CAGJ2AwRWFRERa3AtPwqdBtfVVXFLWYE9I82QlIwh8CbmohKqXJRFiE2n+6pPr2xYPEpUMSKcpvEaH1ePzG69RZ9dMhBDxo0aNCgQTAY0IMGDRo0aNBnP/upnKyqAXUDTdhMZ2sRctasiFjXEKMxmxkCMhFzMJO2nRGCMAqzmkhOKoqmaMYESCgAgYg8zGuGAETofb6qIiJZUs5ZVKAlKNYpMxISTZvpZDZdn05EFUMc7710fabPvLD5qU//+YMPPby20YiAGUhSAwBDMSn+AjEAmmYfaXjJJZe8//0f+NGPfnQ2m5048eITj3/bzN5+w/UFc4HgAwABoE1Z1Yidc8AcgqlJzvP5HMyqqhJVAGBmdy9CCG4TiyZ/vG3blHJJyi0RIUajESJxCJLFVP2JSKjiTAms69pdZpGcJaeU3Lz2vu+6rjc3Npq2jSHMZrPpZJra1MybyeZkOps2TSOS3cK2zmfSDgprO82kV6kd7m4fTF56aKfphLvPL9v+xJ0O1yJmCsXYoo56vGU95vMXDQo4e5FNdYOQaHf37Oz65Y/d9LkjJ9ZnqQMrKxqgIyMQCLkL8CvALjFeLG+qZDKRy8EAAET81Z84/OpIx8QUfUonIoUAZlkEy4gxRDQjY2LzxnnynaOEr2fOeNpmCmRICkCB1UwdHAugcDaf8o0gn89mZqCdB12M1oXFiksn2Cffd/U//sTh12V3E2Ef1S+PLP1sSzeCV1GLMth5uuqieIBuPZotLvbdLrqe9rETy9Mt0P2zMzOX5XUgyWku0jbNvKlHo/HKeKUamcF0OqXOAJ7Pp45MMSd4U+AQQhUlZxEVSYVLxExAAKBQRhr6nR8A+t4XIv9AAVPLKsxMSKricwurqvLPEe+/8SLTzlA5ut3s0wK6vgojQkM1a7MDQHjf3j0zptls2szEDG1h7cPy8EbfLy3A8c185rFNi8/PtPrwO6+/Yl89pixpwiaRqGmlzVmyhAjM7iCjKETDQsQmQkTutllVRZVEoDtD6roKcdGlEeLY+34cty1gjpzKksEAkUOIiChmapCM4ubmxrxtKbw/PzgOs6wDi2PQoEGDBg0aDOhBgwYNGvTW1j33/BaYipLNhUiIQXMrOo+RUJU8l9tai4iAhKiIGRozUU3ZJKOGwJpzTokJmYgJRQwRiEipb7NHAFOxVnPbNv5NnpDYwZqEiMCIgSMZQM5swIAVx7C6wqOV7661X33kmT/9/De+8vB3jp+cmrGYdSOjAKDnIPTxNLzkwIGrrrrq8OHDV19z9XQ6PXHixMmTLyHh6soqEnVTEcEJGG3bcuCA7CbGIoAMEEJAAHZL2kxVswiY1XUNACJCxP5mQ4iej3YIabGnJTMH5hA4BGJ3V5DcSy2UDwBAIslZrWCOHSpNROZYkCwqMktpfX197czafD6fzWbT2axtm5zzTk/pe+DrvVJI+TV+tcXKsf/VuqOM5X++ZD9azKPw/t6XI5SvwoG+aBz/q4/d9L/+0bd8TYTkDryZmgKw4YL/W5KXy8dgi+tuttg+gDuu3f+Rmy893+3pVtWv0rRD0/YH34EbigoAaooFOYCimuScGMHfCzVZVQ1Ry0EwMFMlQoAt1+8bU0sB4l7L95xy3A0A4Gfff80//uu3vl5W/8Ys6RJkHAFk623Alk6eV1jXOR6VbYttTy3v0CsusHXtuz9iYGAiZtaAqWoGAOawlC/eQeNBoZw5s4iYbukO6e8jZiYiPioWAFRVSoK4x+9YFlE1IlEHGpmllHBLILq7P3XVx5fZA+Y3rS1/YYoYcXWVmZipmc8kJ+hd+K1lRENoDbLAXO3I0ZeyQpqn2667/NrL9+X5nKQJYKnNOWVTYS6FCQN0PpOf1swMBpIzAjoj3mzRlGCqIQbvzrGufLGoOSICouOztEw9tK6wSm1KopgBEcSSKvEEVlfDRCAMHvSgQYMGDXqLazCgBw0aNGjQW1T33nuv6kS1VW1YlesQAeeT02ANMQDEkgVmVlHLGpkM0QxUMqKGgKKqJiamkk2VOASmwKySPePljE5m9pZiUck5p5zrmqrIITCDKagREkIgpFhBFp1ICGE0GnO1wit7W6ieevbIfV98+NOf+bNWSYGZWSFrcRq3yNRC5JXVvde9/fpbb7311sOH27Z54oknXjp1Kqc8XlklRDNr3fZF9CFXs9m0Go1DQNWCTShT4zpDwVIiZlVtmia1LQAws5q1bVtVgZm04+0SkdvHMQYRaZqmrgERk5rvh5Rz71mklGazmQM9RBXRQ+IBAFQ1BDYDSQkMRGQymaytr62vr7dt27YppaQqHXDjDe7knVVnN+0WHIHdjbFln6e33C58d/zUHVf9/leef/z4upkSMQKq+f+MEMxtGlHPOFsfPu/yoP0mI2DBBiMg4D/6sRtf9SbZwg1yqwicxdEZ0KpacpOqUq49JBXJ7YXsiQtSk0RFfDKp4wtM1GHeqvLaja373sjK/7dYuZ2NCLBAQn/kloO/9hOHX0eeyPq0XZ5yaWa7scnPJXe/I3q8+1I7FzunQ+n37N37Il75mQupSCuSUitZqtGoqmr330PggssoDSikIJC6PgaAWFUAjozoJuwBun/d/Qp9RrjjIxUEh5h0q0UA8Pm0vUHbly172xp7jDKRk0kIOzrPbkHpqq6YiTiYWQumKqaLU3BpT2AGAwMmfPbk5sbGdHNtbWNz2uRrMW1U1o7YIGcURVCiPgyPUGY3EBIwB1NrmjkBUue8mwERe3EImgaKK63afbQFZgejI1MWySqEmEVSSkzkjTvz+TybhThCipFJiAihgX01rOMYHvqNH3jvL3/5/A//oEGDBg0a9GbQYEAPGjRo0KC3oh566Dem05cADqhOETGOGSSb5dG4JiAisBBiPYpckQFkAdYQQplGqEoMdcWOuwDJQIzMBIYqqGJEAIAqBQ4Q2F1GFQEE85F6HQgW0GBcAShKQpOc2ybNAbmuViPW33nu5ENHnvz9zz7w9UefmucyES7n3M9K2iE7cMklH/rQh6+//vo9e/YeeeSRky+9NJvNQgyEOGsaAPDIs1lxe0WkadqmzRyC28ciklIixMABoDh/2hnT/lX85MmTWURERqMKEXzAVEnDouOna1VtmnlKGZE8fKeqbUo9WjSlNJ/PR3XNIUjOBoZozCGl1Lbt3r17CXE6maQ2zZtmsrk5m898WGIJaL+hELq41QwGAG+7f7mNXPKwto/26hcprsj2lXqSdpcVokf8oH/aIr93nmLCX/uJm3/p//6imRk54cRMxczU2F1IU0GzLNt9PVxEZ7uwoyqA/dSd19x8xd5XsTEuySm3rb93zyoiB1ABA2A2UzDVDAZgKkgEhuDo1tfvv3bbLH6Vi2Y/sAYGCgjo8JTXbcvOQaparMxSW+iqIc4pLqF4u+ri8T//u+/elr39Pmtjnl7HV385vZzRvHy9n7cZvVzrMUhtEtF23lR1Parruq47y9T9ZcpZs4g4UoOJSidPuZn78d31FoFl8OxiKF9/4w2BQwhN04pIfzPvLGwUEet4O9CxpM0s5URETJxzNs8gL4kQ61gxc1XFfRftm8+rzc1Nk2wq3fhYK8Qh6ABLooiw2epjxzYgvDBp9apLRm87uOeS/fv21XHEiE5nIqpibWa5EDbATL2rw1TJ7WdHXYMxsc+wdeBGeU1TW6Sfsau6qRlwYFUTyQg+O6HyT6gQoxhkwKZpN6bzVmWO+w5e/HwzO/TQb/zSe3/5/zzPoz5o0KBBgwa9GTQY0IMGDRo06K2oZrqysvLS2hoi4nhcR8Y8T2jKHAJzVYVxPQoUGBgNqDIyY8JAGAgRjQlCIGQDU01IIXAMIAqaQUi7sW1EjB5/BgQACgEQMQTrqNBIbIRqlnOSZqbtvJ3Nm8k0hJWU2+MnTz3wlcfuffAbX/vmt0+8tC7gA5469EGXL1t+XzfdeNPhWw+/49Z3qOoLx449++yzk+k0xJgli2jTzGOsQmARdeayuwCqlrIQcwjB27GbpiEkR4K6xZBScpe5rmtCnM/nWcTMzAQRVJW5+NfMxMzT6VRVcs5mhkg5lfScdpaoexllaKGIP6SmIo2qEZGqtDlvbm7OZrP5bD6bz3NOItm6KXc9feH7eeacn16VRW79KDLYmvzb8mP33he5Tjc0cesTzi3RuZtuv2b/J9595Wcffn7ZxS7lBSyo712pr526RQEAsY78yz9286vbEhchLcKVDABo2LXPOwHcuqF5CM6uFREk3GZ1fT+V1ZiDmaoYkJcjEJEAAe3lixNvDG2vXiyfXMWIRgD49b/9fZ06uKvW53krA9pw65b3EIVXkL0sonmHeqjKWVf3ii+4IxB9XqAOkawqkgnMCCDE0J1UDjtWMyVEDkFUAUyzGHb3jo7XVDzVMlzWCw+LwbPQLeSQjWVjernq0N8H+oh0/2tJRiP1T0TAbdUXAxAVRCBijxLX9SinVlJSyP2y5c7f3QEFbK6WZvk7L5xpcj5zaA8HftvbruJxrAMEE1EBwLoaeRuNx/dN1c8WVUF0U76c7cTs1eGcs4oiIUDHHOk/fBeIEY91G5dhjExIVVWBGRGLZlINKzUirE/mKPrSC1ceOHTolKx/6lM/87M/+9vnfpwHDRo0aNCgN4cGA3rQoEGDBr3ldM89v5/yvDl5EDiPR1UkBZmvjoMJquRRXe1ZXdm7b1+et5okMFfEEdE0oymjDzUyA1VR0aSSgymZgoiP6xIpQNJQExOCGoACIBIBoolozqCKiDiqjLDZ3JhPNuezzTSfpjal1pj5pTPzL/zlN/7kvq8/8JXH22JJljRZ38Lch8vcI2bmD37oQ+977/vM7KGHHvra17+Wc15ZXV1dXdncnGxubk4mm/v2XbS6ulrXtUiez+cAwMxOgqaucdu/bItmFTGzGGOMMaXUB+uouOpARAWdgRhC8FmCnvCeTKaeiauqymNxvoV1jCLStC0AxBhHdd2mpKoVsyOmm6aNMYxGo5xz0zTT6XQ69WGDoirWxeFKKK5go/F7C2X+XqgHh+zGl97dBdseVCwN/dCXIswMXi4a/2r0jz5+y31PnNycJ3ea3UMlJkfKqHoNZUcCujTOAy7Mcf7Fj95wcG99IRsTqhjrGgDQsTZmWcSx5VJQrKX9X1VjCGbWNEYUQn1Br3thwlBFFTHLZb/1ydBdOblvJC3xd7tIuxYjt69+feLdh+687pLXZ/uWNGll+TzcdjswXRjpr9AQgNuN0V21jJk5m2N8bgn3ZQ/aOlv7lTeh3xQzA53PRHIGxBADMSOiqpkqIIYQR3Wds+ScU0rmr4gOk6DuUOYQ2Es1OWezAkrqWlu8ioNEwBxUNSUvXrKq+LvsicnM7Jehr6HPWTOzt9eMRiPPU2/ZU2ZooGpmYiYAOB6PWsTWIGfHcQD4h2gIKgJmiCRayNYvrs/WJrONzTOrq6Nbbw11CwywwiQqpkqYCBHUkIgAgZmIzbRJWSELgKmKqqogF+WcVSUw9970wo43ACyA7KZplj36xS61NmtWk1CNag6rFW/MQUFOvnB8/R01r+fBgx40aNCgQW9BDQb0oEGDBg16a+mP//gPzKRJo8hpdaWuUE0TqFhSVGVQyqKzeauac9KcGpE5AiOASGCuQkQCA1UQHz9EhM6ZJPS2YAUT9C/roKBJu3FjSOT4i5wSIq6Mx9JsNilNNzaadi4qe1ZWqoonc/3iQ9968MuPfe3I0WeOnWwMtBgUffxZALjEZJGqWF166aU33nTjnXfcORqNnn766eeff35tfe2SSy4xsxBDVdcxxn379uaciTiEEDisjFcuumi/Z8GC5+MQPcLsvjaYubtRVdXqysrm5mZKiUNgZuyGE4YQsiQACIFVS0+3D7MKIQJACKGqKjOo4pw6SmabEocQY/TE3XhlhYk4hJSatm3GY805zWbzkydPbmxstPO5TzX0r/+I1PFd3Q7o8MI7dG5BwnNxAHFp/tTSo27cLP2+y1px50P9MzwRCIiEO/AF2wfUdZFeUyUvY1gZJLkwMZGLMU9EpT5hS379q9HBvaNf/OEb/s1/fAx8IhktooLYNdFbF0tceodaBmt2KdorLl75ex+45lVvhouQ+upITknNVNR8nOcSKJuIQgg5C4BVVSSiQOcC//2eSIs/CLTg7pREJW6fxPaGU3cTK77z4oTszk1C/Ac/fP3rsm3btD5LW53lc/X2ty1nu4F9zupZdwexe55tQevsiN777LrdVtMB9z2FfQ5n7I7ViMhkc4NDCDGO6lGMkasoagCQJSNhVYVYBXM0EBQaRbFVOXR1Tezhz14+9PGGMUanUhQGMlPnO5P3uMQYc845526YIRZbGbGqqh7T4ZyKbQZ02Yje4lVgIgSMMY5Xxk3bzGezZj53419ES+nNSpeFmCGYGJxcyw998/kza/e+/9Zrb3nbgUv3VJBnpO1Fe1dBNTc5dMo5S84iikQI2LaNSMfEQSREAyCEEGNXkjARzZKpmMwEAGqa2gQAzFxQJOSDIiynJJoVNaQMFAipJpCMorhyZDp9x8rk6N677rrrrrvueuUDPWjQoEGDBr1ZNBjQgwYNGjToLaTPfe73VBWRVduqCozQzCeoCUERAA0ILGnG1Op8BiBmGSQLAgOgKYTIVgOagoqJfwtmo/LFlQnMVIUZqRgJWbOIug0FRCQikhoVJSLTYGYgGQMHq9msGu1dW58/9p3n7v/ytz7/4JGjL5yZteIdy8tug3sc/sV4z56Vgwcvu+2222655ZabbrzpqaeeeuGFF46fOB5C2LNnj5uVgOUbMvi3d4DAEQBUNYt4us0zgk5zVtUYo4rmlJi5inE8HptZytmTp55iY+a6im1KABYCd4wO7A1oRIwxumnIHLAbyehOXG9D+PgmZs45ORtkMpmur6+dPn1qOpnu8GtwyYjvH9lu5Z0PdeLcPOhtvy9s33N8kW65zsorfe8ASNgZ0P0yuxhQSF2skwkRQcEzg8ubhAAISFyMTkSvL1yQzflzH7jm01899typKTECEmDpZIfOgFZbxLWxa0WHLkrv//xvPnbjKF4wBwN7gYiAmr86dSPC+oGEBc+C4AMtX0dpNxGuKxt4HLeL0HaHb22WzkzbaSuilrN2Z3RJuHcACbSu9nLHtecROl6fpae+O4EFPWCLfH8yYhUoMq1UvGcUVqoA/Tm7/VpaXH0fOXz5tQdWz2N3dDq50XzjubUnX9x8/sx0Y5Ym88SEq6O4ZxQO7q2vPbB69YHVtx9c9c04p/c4TVu307beMBe3i20Wsy3Ril9eOzkbZyFv7FaIWnrerneMLQ8jntP9C7cnrFVVW5EsIupheyxVD78SAYmYSA26wZ0G1hGdwJPL6J9TAMG95hijLxG6CQGLO1nnmLtV3V9r5SUXBA/15hi/ELxCiV2x07oBhojYzb5VP0KEiARgxiGYgYhKSr2/j4DmNzwjAxGAZLDZ2NET6y+dWoek7aw9fO3BEbU1tghKptLmKsbAgZnaNolImTqI1LZNMcRxKYyO6EyqRWuFny2lHQTMTEURUclJU8gheKNSlqSmgOAetyGBMZgoBtU4fliPhGsO2YvncJgHDRo0aNCgN48GA3rQoEGDBr1VdM8996i1RElVOXDObTOZam7QEplSSW0ZAwSyyFgFCoECWSCKTGAUmJjdpyVVCyEQI6gwU2SikvnSUNeIaKkFUzNBVPDv/wCBgerIRIiECDGOxhfV++qRJdFZ2wo/8+gjv/W7n/nykWPPHFvLpuIAjw7WueiFt/Jd+ODBy37gB37g4x//eFVVR44cefqpp8+cOXPxRRd7vnJUj9S0zYmIO36uAECI0cwsZ8vZnLzBTMW1VI8q55SbpvHw2rxp/PVS21o3kNAxsMw+t1Ddeg4huOmsOnNzIaWESKPRCACsM+OqGHsbom3bpmmQaGNjfW3tzGSyubGxsbm5Kc6PfoPHRF+1FhwDKLUM7GwoBCwh5i3yHY89inSnS4XYuz8AAASEtBORcV6KTL/2iVv+6W9/gxBtgX4G6G0jABXxmD8BEBJ7Jaaz9t75tos/9o7LLmQbXGbGPjKMSERzl4snouAkcSzhYkc/u0Qknw+V5NlT068+c7p/k76voYQ0vZrj3pMux74R0SeUjiveOwr7V6srLhr5I5qFmKjjD2iWvvaQsvyHB57+9/c9dXraIiERmYFkKc6dChIhkqoCAXFQKVfrQ//ib537O/rWsbVf+fdfNlOT7NtKMZqq5QxmQATsdjMioYqY6rgKN1y+79Rmq8WkI4dDWHf4/dL+yduvOo89C2AAf/7oi//h/qe+9sypECKS8xkMDDiU+kQ/XpUQb7x8z37BeD0AACAASURBVB3X7P/wTQdvv3Z/ddbTeL3Ji1dxR1XLz8uPn9fWblnfTvrNjsLYLu7+eb3Mzh6JVyU1tZSmqm1KsW337t0bKjdwRSTRkgHNREzsez53nSsiZcysqvrHFDGDl3NiQECHcgAAEfm1RoxeSnTHtsPMFAPaf+jHFS4tySI5ZwGAGCMzOVCKCL2QRESaE4BVVeVNMHMRyeUcNnTzmwCVANUgmTFjo5Bn+tA3j25uzFdWVw7tr6GKzZnNiFo7lkfnPpnADEyRmYnJ7ySIEKqK/faSRVXmXf9NXVd1Parqum0ap1H5m4wxqlnb5qZpAaCqKxU1MyREIiT08YVqOhMTGgFTEgOmO+2RdVz53X/5d3/6n/3eBR3vQYMGDRo06K+OBgN60KBBgwa9JXT//Z+azWY5jzXCeCWCCSsLG0pEVEIjYkJAhAAWCWOgOnBgCmgBISAQGgMQAhIaYo2AgT2NSYTEhGbQDX0C9SAXEBKyW9YEzEAEACiCZhYiAlrOqvPTa5MXjp388tce/+KXj3zlkedfPDVpRa0EZKHrNSZbONG2Z8/e295x27ve/a6bb7752PPHjp84/uSTT85mM8nSNI15gIuDgolK3/5fEtChCiEg4mRzU1SZ2Ue8MQcRMVMiyimntp3PZo7LyClJZx9jN5ZwNpupidOZoUAw2TPO3o4tkj2Ya1Yg0aaaUmpTKsHnEObzedM086aZTSfz+axtm6ZpcspdxO5VH/NdDNpzedo2y3u7z3SWsOT2WDTuQgdZkBdwhyOG/avthHL0sFnrOaQ7Zaaeee5oAH1T+4XoQzcceN+1Fz3w7ZO2FM3EzisHgH42oOSsZhCjG15epfivf/T616SGkFPbNI1XbsBBFmpmJuC21GJ7XKY6zxkQLVbn/iqPHlv/n/7wSOcto5kRISFmUU9YF38NPDsJKWcEICbsZqz55jHS1ZeuHLp4HGKALnjLRBCAOkbK//YnT8yTEGAIgQjVrFRomADB1B07QhUvLRDGV2FPIiIHBiNgtq5ygUQYI6LbZJ5FLTPlDLFVePT4BhU/Ed2XXGYmIOIo8gdvPHDum3Fyo/nvP/W1bzy35rcmkQyCPd5GRLYh0dX00efXHj22/lsPPLNSh795+5U/dcfbbr5i7841i9q0XRjQiAjmydwtYeezsDXOfo30mPUljs4Ot3nHCsx2e3TXTPQuy+xSfTrLFm55soGBiYgBeIq5ShUzc2C3jE3Ng8YCnlxmAMyqfqC94NEbrJiSihoYpcTkaOkSW/YGCL/MAcDT0/0Npzeg+6Ogqr4ry7XA3DStSOF7xBjLBd0Rq6hY1RBDyKJAXK+sppRSSlBoGeWM8fIuAiQ1BQsEp1r59otnqi8/eut1B2+++tLrr3zbakTOzagKgcjR2AAgWUrhBcBAzSxWFQKmlFNOKkqEnsoOIYQYqhjnbZNyVlMEJOYqVmqaU+4sbL9kyW+VZqBmRMhEew0zhLnYKOu0VVUbVxtR8LN3/cwn7hpg0IMGDRo06C2hwYAeNGjQoEFvfn3mM5+ZTefjlXZjQ+q6ruuYGqGAIYwIlMiIkAITISMwQECMTBVTJAoIZMqmkQBMTIUYkQiYjNAAgAQ8v4aKBmggKWtKKhIYibE0CxMCkwI6NAABFEHblOd5lvQ7Tx176OuP3fMnD37j0WdfOuOdxqhmhECFNewJO/+qzRdffNE111zzvve977rrrhuvjL/6la9+5zvfOXPmTD2qQwiz+azPmqmDkztTUkTNjJBH43FVVbPZLKUEAArAgUejkYh6FzcYYGdoOt/TVKmLLTslVFVEskgWKX3W0JESACDn1DRNjJWZzWZNXddVVZlqyjmlRJ2TPZvNJtPpxsZGTq1IdoPELZ4LMC7tVRvQO5+zcF3P1qqPu6x/x/JnWcMWF2yn31TMHUWjrm9+B8EWwFQRAc2HgKmJdlyKC9KvfvyWLz7xYsrWB7ehi4aCQazi4nwTQSIANDVV/fF3XvGut1104RsAACqaO6N5ucffzLIYdQFL6JgAZiop03lSOHwfQgexBTNEJiIGECxcbVpi2hSiBgBx2ScA4BnSZ16aPnlyMxCbmZgyIjIhk1OrzWOnAQiICQkpSfaTiJiIWE27yGihKXS0hPM9jRG7nWNgqpZFAIFC8J3mq/MbBS4n6A049MTbZADYIa0B4I7rLonnHK4/sTb/B//2gZc2m1KBYZIsBRDDCIAm2p/SfWeA71BEnDb5d7707O9+6dkP3XTpL330xsOH9i2vfNLk3fzf7Q8tn7c7t/Asy8MOF9t2vb1sfaBnB29b647lzvlGde7XsZmBSTYVAbCcUoxxNB5544t/FomKFkC8AmCSUlz0G3s/exAAlh1nT0b7i3RRaOsbEaDQTrS7AF1KRAaQs3gsWFQBkKlwMPwl/Aczk57L4SBmIgAUA+IQqppCUptpzqbSgUtK5wgiZjNFM4IkcGx9Nn3s6KxpKdRXX3f96KJxrU3NxgiE3vCDIgLlgi0NCn3K21PSpbRW7Hggxjgaiak35njJ1ottAGimIhJCJGYDy6pZVLIEprquwKhVmLa5yQCTjWmTq0zRcJ71U//0Z372fx486EGDBg0a9ObXYEAPGjRo0KA3uT7zmc+ANk07grwZohKYtFPUhGiIhYyBHnAmCISkBqopt0ZkxBQjqIBlIjTLmjMzIhMSZUkiGQxUs6qwu7MIs+lUJMfIWFdILN5nbgqIbdtONjfGo5XAoRVpkk0bObU+//wDX/+9T//Z89+drE2yUQBVBMMOF0tEYKDm3/M5xvihD37ogx/84Hg8fvrpp7/5yDfX19fbpq3rmpDAAAmrqmLmyWTiDjIAeEIT0USkTQkACLGqazWbbG5mlRBjVVX+LXo2mxFgDMHJJD48imMExKZpZrNZj3JumpmqEPFoNKrrygw8+0yERDQajaqqVtWUsoOejYhDGI/HIYS2adbW1yeTyWQyaedzNTFT0N6KYkCA18I/fYNrZxTaRHexqj1Qh9anCHcuoCoIhj41TtVMTeXCt/DqAyt//wff/v9+4SkvZjimVlVMTQtsAxCRmLUgvymGSGb/7Y/fcuGv7qqqGGOEzk8FAD9XTRXIra3OL1OlwERMSGWDz1mIUKAl5SQ0QsIQSteCmeasAGCA6HQcLalPMwMQ8SSpKooCKJhYuRY8Pc3ExIxd/t3UvKxkhKiIiMzEzEhMPsgRi0Pp8dXtMe9zkJmmNhFRjKE84JPeHLa7AIyYirhRbZ797u1mJCTu+i+87Aa3X7v/3Lfh13/366emrZ85HvBFIgBTVepMbhVV1Z5gXlAGvWusZghfePy7X3j8uz/3wWv/yx+9aaUq1I6Ned52BdkuiIzFVbZrEWinPb3r8p39uh2A480uW7eh/GX7hsHWs9F2Hs9dNv68ZV6lwtQ2knNKMUuuR6PRaBxCKROqihlUVTQAbROR11kAup6GZYaG29AeqfZltISmKQSnMAkzh8Ai4u+qnFSljOJwHmbmpmnc2/XPCwDwmoxvNXkfABaIjp8bbGZmpYfGrJk3OTn52atEoGAGCoSGlEzBQA10Dt946qXJHC85cGl8x3XXHzo4Xz+ZZ1NTqSPXMVaxMijo6Sw5talpmxDCqB6FGNyI94swtY1IbpOMxuM6jhTMVM0sZ3UQBxH3XjwAELMakCkgR451qFPOEW3vqIZZXgkVZtlscIYppVjFfPddP/mTd919oQd90KBBgwYNemNrMKAHDRo0aNCbWXfffbdpg1RTfgkCjLjGPFXNgYxAfSgYMGIgUkYCA8giIIpmiJSIgCkSBnS3K0lqYxWICRBzbrNkgDIj0JAEAQFMMoKZQZtFwE0jAgDJklP2DmhByBlnjR4/uXnfXz78hQe/+eSzL80Fk6KCdhTYEo+zLv+6umf10KErb731tnfedtuevXtfeOGF5184dvrMmaqqLlpZqaqqbVtVdRAzEQGCu0zuFxOWR1LKHEIVIyDGEJjISgJ6bKYSq7qqmchHMLkPwd0QKkIMvjZmZ/KquvUQEMndDfcm3I+PMahaXdcxVjGGzpXQppltbk7W1s7MZtO2aUQFOiOvHDzbzZt5GWvm3AybnSvckVDezd1z7C8ut8Yve1jb/Kx+sXP2CZeBD57hQ2JYwIcBAJgJEBXMLUkPm+/MVzJxP6wPCM0KGuLC9QsfueGzj7z40maDbhEamJG7MNBtffCZk1mIKDD9J++/+tDF49fk1QHA+c9lWmY3zLF4ZG5UlhGI7mZZAa8vmCfnpHIsCvQGCNBUJbWqZlroNOBHBdHd7RLAJAIzJ8m7cYxmaGamoAQenFUwcF4NmpWLWyUDohKbuY2mVoKZ3gWAZgrm8BwrKz8/FWqzc3jLGaNmHXocewqBmY91LNPfVBQUzBBQVawbpuqm5LUHVs7x5b9+9PTDR091KAs0ANAFisa0O37lV4WOkb1dhT1jv/XA01968qV/9ffuuGr/CgBszlN5n9Bfed4DUH7e8nz/qSuZnC34vJvO1sGw29I7Hqbt5vIuUA5zUj9sX+68XOlydpmWyqVpaVYZjUZVVTERAkjB94N/+JkWsrnXA/zkMABA88+O7m31XQilWlO6HxYYaIQuIk1MVoBURoQGhoRoPt+vz1YHnyXQl3J6s7uH2pdPMUQEjCGmtk1Nk3NWzd2doNtHWvZUY3B6lp48cfpPv/To+sbmSzdesS9a1CbPNldHcXVU1VVtKqpKzFnUOc4cwmg0ImYEcAOakHJOqqJmzbzx4paq5CwimZCYg1+ZXiVS853hpTHKzO2U/b6FxJa1MuMqaG6mrYUqA+fTdsldd9111113nc8hHjRo0KBBg/6KaTCgBw0aNGjQm1b33PPvRKYiK1FOB9ZRYGgmBolAit+iaioYCJiByQDUVHIGNSYUJEDIZlZFDJwkS2pzSpYjBwbCnJNoBoDAIQQ2VQXwoBYxG6KY5axcVVyw0AYc6tEKh9ogKNraZOM7R0/ec+9fHnn8+c0WkAkQUs4LpwERENWMiEZVOHToyne/5/aPf/zjOecTJ048/u0nTp06NV5Z2bdv73i8UlXVxsZGSm2MlX8T5sDuHxEWxzjEiERZ1LpUWxXjeDz21vve//WlvUnZv0m7v5ZFQghuEjEREY3GtZYsWPb3vrTtJc5pZisrYzfBRSSl1LbN+vra2tr6+vqa5Gym4Pb/kum8xYw+q87RmCnd891vnY35inYeLoGb+1fEDgaMAGilL9+6l3lZ8sbLGVjEnvosG8iEBtj5M+WIuK9phSbsPN+t8/V6J7uQFRBxAWi+QK1U/Ct/7eZ/cfcRjyYWu5wIEbOImiFAYA4hCGQA279a/fyHrnlNXrrIbVI1FbVCaXAD3LgzrjyFTUSSk4NckM/fr+1NS0QEUBX10LMZqFKIiKiibtualR1dEsq9N+eoWbEOzWIOB9GsHT2gmGuSExgAMyKBue1rqASmnUFMTrvpV32euw2YSdUki+eLHbsAWhxtQKLgW4mmBqYUyK1xVQBSAFTJpgUr7KMLr7x4dI4b8NVnTnWFAmIv+qkRExCgovbYawDw2hUgUs+73yEDBPjO8Y1f/LcP/u+/8L7rL9szaTJ2Vx4uYM39FVfW3F8s1jVV7N5GsPMFd4lC71LUeJkN3rpcV8g6+wuC6ba7mh/6Hcvtsq07X9oMzMlKKTVNoyLkPA1EIzJzIAarlcg5IyGhiYHPn8TecgbDEoXGUuxBr4QpKiv7h0Vd1/21gIixijnlnDP03QlIxBRCmTfgCWLm8nTfZlUtmKbSvtN50CEEDqO6TqmdhzCbTdtGvIkAEMz5O+qbCmLQIHx3Ov+LLz9+4viJ489ffvuNVx1cDTI73Yx4XofaP7VViaOqpVxg6yFGZEI/URctFIiIbduYWV2PREQka7HsSSQTc13V/qHZNHNEYo4xBDPLIjEEDszECkRISLQaELJM1AjCk/z2q+D4K50YgwYNGjRo0F9tDQb0oEGDBg16c+qee/6dGTI3iOJEgqada5qgCaIiWPSGXoScsqSUHNCKGIiIiRHA/Auz5IyBfIYehRiYOUaOVSXZEZbqI56AGJiBGU2BCGJ0MwCZNCdt23pEGitNwmHUCk2n088/8PAf3vP5bz91ctKYIKEjFgBgq7lgZvsvueT6G278wAc+cMUVh44ePXr8+PGTJ0+2bVvX9Wg0ijGKyObmpoiYwXw+BwD0+DMAGjCzz0qKVQwhGpLk7CxmJqrrWs1EJKcUqyow55yhYz27YyU5q0hKqbicZj5xblRXFKg3C0JgZq6qSFQguZ73XF3dk3Oez+ebm5vr6+sbmxvNvGmbRnIq0bDzDPi9kna6PK+QfX71oq3DB8/T8PTiQFkTqwIBAPoJiItO/5JM5EWwEzrQ6tLKPJhbzNlCoX3t3uiPveOy3//Kcw8/twYA1k0VCxwK+RWgbdvUJgJAhF/4wQUk4TVRlmyFt7yw8Yrf6zZZwQ6AGRKRdYxmrxKdo7ww46t2OAYSM7G/X4NcKMm+XAYVJSbPS8LWcxgJGdmMzIPYxIhgqkbshiwyu2/9/7P35kG2XVeZ5xr2PufezDdY8+RBtiVZlgchz4CLsYxtuqCgaIiqHiqK7miqqruBJqKHgKjoVkd0F1ERRBFEdTcBTRRFdVVQIcAFGGxkC2Rjg0cNz4Nk2Zpn6b2nl+9l3pv3nL3XWv3H2vvcmy/zSZnPsrEc57MtZ94894z7nKv7W9/+VrmWjkqNAbzqEQDAwBDIzKyOswNb2ldyPEo1hYgBELmcLy2m8hKOUQob5lEhxQNLjORdWt2HbEem+23teHKWkAjUDFSyOPJ20MyBdSX9mZgQ2SuDhWyqnrW2gQJvzPv/9nc+99v/zbs2F+X6uoG7LFSHvZWkY9uxBlxi6P3rnEz8JaAScAEii+1tVZ1OJtO1tbW1qWdH5CSIBAhepWBiKeZgbZrGC4eGJQLeI5IHe7IHwVtr/quzZv+r37BUJ9MwcxmASN7ZEgBCYET0B5fWPrer5ZxiJ65Em5lSSjHE6YXTuBm3NrHbVkXvOykAAIFKdgyaAJhBD/DEyTnqsxddePHFF1/0mle9YrHxbJ6fkayBMUROORPx2tpExNQADCRlEVERd143TQMAXj0FAKKeOcTYeOxGztk/Z03E7ylCZObIjAhqRmCqmQSQGE3IMhiREogGNmR8J9x9Bo/86c0/+Z+MDQlHjRo1atS3r0YAPWrUqFGjvg11663/VoEJxSwSUYiNpHnuMwAGZkAGMGwaDjEwmiqYMmFkjhwIgBEZHbUYmLYhNE30RU0Fg+chBxYxVTMhUEIAZogBYgOSwBSYPB/XVNCUCczIgM3i6W154qkTd9z91Y//9bEv3PPQdiYxMgCtlkerNmQAiDFeccUVV1/96muuu25tbf3UqecefviRjY2NxWJRZycTAHhws//u0+1FPAmBI4eUU855e3t7KtOmNSBKfUopmRk3DRHlvs8piWqDSMzS9yoCiE3ThBAAUUQkZ1V1I7OZiVlKiZmYCxozMxFdOoPBXwQzTSnN5/MzZ85sbJza3NyczWYq6vP6B5j69SHoFyTOe76yvzUNDQaXDkgsLsi9TJHDwe+HWGGlZQXEFwN1/XnnzjzfmgusVjA0RCI0K7bAF0sI8PPvufanf+vThgiA7v5TLKMW1FTVTYPXXHr4/W+6/EXbMAAAqIiKWgWgbqTFavoGA0/HLmk1qgCGSCtt8/anEuZcPKdLwzxRjUtWMDRTXFpD6/4sN2RuxwREsHJDONktCSJeHTJDAywr9s0goj+RAAgLcC/cuY7AA1u6ff9xNYEGlzbvUufwiRKDhRYBoRo/y41ZbLAEBmYy3Xd14fAkIhKggJWpAzXkpPxS7NGlAyKZGajsx5t8atb/4i13v+eNVwyvDAHOO2/jMkLrwb/Ixa4XX27pXZGh4c59Pr8j8EdxiYdAAKa2adDrAQRgIJrdBwxevBFBBCIWFQMzMCLMeQeA1jpVJYRARB4DVS5rvQx15NenGiIheYPUnLM/6CpnVi7VDj9MG6I5wMEuUUrlLYDIMYbcZk06fJS4D7qOBQXIAKcXyU5uHXvwmcl0esEFF6wfumhtuo79LKAgWhSlEJpmUg7S3BjtDREVACdtC4ilPS8AU+ASXVU68eLqLWVgZsTMxD5JQ0sQPyJh8OlXYJJl2oZpy71AD3QobwOMYdCjRo0aNerbWSOAHjVq1KhR3266/fbfToIkkmEd2EIIOfdKBG3L6GkZSIht0zQxMhMBEEJkamPThpj6DlUjcWBiQiKITIG5GKw0Q9MCIYgQAICCZMgd5B7QgAnaCL1AytD3knJOWVRC4NjEpCbKnTWPPP3UJ//62L/+Nx946vjpXhEjo+Pn6gT0r7EeXjGdTt/xjne87vrXX3DhRZ/85CcfeOCBlNLRo0en08nW1pZ/2z906LCInD59OoTQNM1kMvFWgTHGtenapGn71Pd933VdjDFaAzWlcjqdTiaTtm3d2tw2jbcHTCl1IlpbKoHb0PxLde0E5TOmt7fnIYS2bVVzztlzZqHSc/855zyfzzc2NjY2Tm1ubpV4hMGSCQCe/Xr+Zt09Ui/2kO1jGYRd5AuHVA2rOBeH5A3EYcV4fkyoxAV7KIpz5+JfPuugVhIDdoVvLANLzMAQ0cAbV+qLa9u89rLDf/emqz5wx2OlsxiAiCD7hAFzaGSqP/ue65hePOu1S02yDNEpZmaiFAISqmgFvmSIYCA5gRnHWLNSDiA//+XKmnqUB8cGAby2Y9W/TEROafXsTo+4ZKClHoOmYqoq4lZiNSUBv+ol/ZyKW9kHQ7nSqogKULsWwoorfp+ykrDsHU3NPIq6FiywWr09+ELNhzMOKSu+YM1+BkMwM8lh39f30qPTIdKEPKKntvIbUkZMDRmH+tn+D+7eJ8/c++SZXYe8R4UG6UBh4CtvXNaHDrD8879l9SFz9mI1UGKHDF4cAg1oqlk1p37RLeJ8e2069d6eUCqIOaVSvMTSUJQJS/Z6Le54OAsQIRNJAccWmJlZVP2jYcjNIEIf8EO+M9bIGhGRLDGGEIOqiqiqlAjyldNCRIjkdxnBMp4lBGakZjKFDvu8DT4mZcepMQAB6BE2JX/y2AMbm9tt27z7O1535WUvSxtPaz8D6YEDxRhiwxyGBqG+7zmllFPTNFAN2qu7hmhISLVPo+NpP2Zf0D9DEVFUc0p938emYeacMwOsEVvA7T6dWQhI7i0jwx/9ix/9u//LH5/f1R01atSoUaO+lTUC6FGjRo0a9W2lW265ZXs7T6fdAtYDamibhoMpgHII0yYgIjAiE4KZm52JiImInKtkn3OPRIbeqQtMRURjDGCas1iaEWIkSn2fU6fSExgREIP0293GSU295qTegBApxKgScpZe+ZGnjt/1pQc/c+f9x7704DMb805JgTSrI6jdeOTaa6994xvfeM0115w+vfGpT3/m5MmTfd+HEPq+Nw+GnpQkVjOLMTITAOScVDUEbtvWTM9snjEzFXV7WhbxpogAMN/eXnQdIS4WCxEh5u3Fwn9VVUD0bA2rEc/e27BEOfd91/fugPa3uz/af/AwaDfcbW8vtrY2F4tF33UF1a0GJZdv8zt49IstfN6VH3wyfl1ZNeQCrFiYBz4x/PB8dk4rznFTdUuvIYLa4A/1zGXx4eSmVDPnO7QCAQv7Nau7pSUs5cU+oz/z/df++Vee3eqcw4KZoc+OZ0IFMPiuay9526svepG3CrXKUBH84LPHEpkNfl4AbHk3qZV7e/8bQbd/GqgpSKkGOIYGQ+/9aAAmQ2y6ia4mRSB5bvtw5hEG5FvKC/6fAvSGka8iK/nToDmXmRDMSCVU2lRM04FO22DNrsbfvThmOcx6D5rakNxhZhWvu3nV39JlPbS/HXjLK4+CqV+rcvGouryHGwnMREXBzPM00FneeWtgiDteOYv0HgR2Px8yPqBe0Nx9oCkUB5cBgA+ntNie5RSbdjKdtm1DxCkhM/sNbWo558lkQkwpZUAgJmZOKfvHEFKtrsBwO4Ko+KnmwGCQckb0+Jji5IeaE2TL0YV15BeXtKllyX7nes2GiWOMiAiqKWVn3szsDUd9Fk5KnUre3TnAALKBKQSDh57d+OO//MJ8kd51wytfe9mRpgHta6qNaUq9qqmUJBAvtQJA13X+LwZMpAAp9V4CdBd4mRUE5k2JiahhVitdFsgbM9ZHhAGU/oqIQCSE0+mayDxnaTIuGuAz+qGfff8P/6sPfwMu/ahRo0aNGvU3qRFAjxo1atSobx/dfvvts9mZrS1gDkTQtIFRCRKxIUEM1AQCMEZgIk3ZVECsdCBUUIBkSGhAKErqeMiAwJjQJJhKSj2ZMhGF2M1nfbdAVGbkQCiacrdYzEWyaDZTphBCRCIAzmInzszu+cojf3bbp+/84iOPPnlSwSe9o6gaGCI4UPRvvJPJ9Kqrrrzhhje8/vU3qMqJ4yceffSREKKHPvsXdU/nNIOUEiKura05uHD+625od10xMSI2sVFTyQLoX91JzXJKqup8Wc0kZzemIVEIwT1p6s7NEqqrWWTAzf7N39tJOaceIjtFpO+7+Xw+n89ns5lWhFqMl4MQXqSs4udZwwr+2KE9+c4uB/SORc+BdN2BjLh6JANIWvnh7PUP/kozwNo5cEnl3FjtiQ3VZG11W1BiHVYSkc0Dh8vfkV58on90Gv/J91/7L2/9qppCsdUqAiMhEDHQf/eD173Y2wTw6esDcPdIAsJqT3cEZm6ydAe+L0qIhAeLonbbpmopIJnnqJsiEjEXPqvmlQGoIRkrrNAvKKyAsGWDyururMANAXQlEsIXc/ukt/uriTaO+QxgN197AbnJ2k+R57Kc3eAOa7J2OX4zjxDZgUEHxGgAhNSls9OZz6VXXrT+ple87IuPnS427CVoXDrF/aYyNTWt9thhOsA517wXyK32e5wR7AAAIABJREFUVSphLENIy54wd5VB79/pvCe53o2V95Mistd2d5r2/dLscR72PQzO8cwzM029pKQibuWPsSHE0DTMDICqmlNoJy0Rkg8f5iZG5gRgTWyISf0M11wV88KNNzNkVjW/Z2srv2ECB6xOEVCvvZWtIBioKgtzYETMKQEAIjVNQ4imikgqUsp9CAAQrfXzlwFEM5THwDKQxW/HEMLGdn/3/U9MGjbNTbz2ojWaYEBJwQPdDbJoTtkAiDCEyMyIlFICMCb21g45JQNFACVEJMk5xFhmC5iqgZCYqpvBgdkfB4TIHNQUandHQzQ1I5i07SLpXCBuZTgjuK633/x933/zx/Z7iUeNGjVq1KiXgkYAPWrUqFGjvk108803P/30Y5df/grE4wrWMpEm0Oy5tAiW0QwNwbzZoAMPkUxEQhQItcAeIwACpz0GajFwIOpNRLKKTNoWQuwkLbpZzmltbcqMBtr1C5EEhIgYIBBi20wCx65XwMagefDhxz57x9du/+Q9sy4JoCGWoAVwgyMwMQCIChhcfPHFP/zDf+eyyy5Lfbrr7rvObG6++tWvcdMrEYtkEXV/Vs4559w0zdraGoBj39ISMOesIiGEJjpTKNkChuSUBxFV1X3fVpssSc7E3DRN27bMDGaiWnzizCXzMmdmjk1DBGbq4Rsi6tmg7tidzWZd189m88X2toq68e4cvb/OSWp2Q5w90E81x66uZw8/OdJeMGYX+96ryZuVkAJET95Y3euCe+uuOBR1OFkZHVLl1iuW5dVXCAlCCV1BxMAkaiJSNgtAzFCCTdCATAQKJ7WS38CECASF4riJr1qEX2T9yI1XfvDup7769BkwRVMwBDQ/Lz/xtpe/8qK1F32L4NPwPZ7A+57VnxGpYE3E6otmAHeUixsZD7ip0hbSzJCICc3ImTFzBCiMqRJhZA7AXoOpZaQVpFiKAkOMMpGpIZjfyYAIkAdM6odjuJK44BMywCEkEgegg/7be6HOyARAAGYgy6znelObmblP2SrvxoHha9139iMCoufm/ZUXTPe5B7/w3ht+5rc/65G6oGWltRBlbvN3fkfGiEhMw11+rhQZpD2QLwCU9TOpKtR2kp7TsueK9jVNYffWz42bX3CFZ+3G2YsZgJVHkH8erYSv2M7l9titXa/YHkuuuNoBLKd+63RazOdN2x46dKhtmradeM0BAd3R3LSxdAhECISRiRmZCZBSylkyVTc01aqX3xGlFWHZYyuTabSMKERyyuwDwOtrkktsBRMTkRuxfVpPre2UskzJ/lAgoul0ysyLLi4Wc5NcGhKWs1hM32tra2i2ubl59/1PzuYLJH3Tay5/1cWHqVtESxEthKhmfd/5HR5j0zRtDBFBc85d2p5MJsQMpgAGaComtVVjCDEw52ySs6RcTkLOQqRSM6ANI0d/vIipqCKzKYjCtIl96jNgPhqPhDPzHPe4vqNGjRo1atRLWSOAHjVq1KhR3w66+eabL7zw0H33PXjBBQ2iMYZABNaRJgQjN/SJqCmhqTdBIkAAMiOAgBipcCMkZHQi7OGV4LmnaIRNA0iRiIiRcA2nam3TRvds8SQoKIAZGqKBWgAmY2741JnFo48/9ecfv+vTn793c77IRgZkgIalXRICGKCoMPNkMr3hDW943fWvP3LkyKlTp06cOJGzNG3btu2QhkFUgLBDgel0Wh1nHnZd8FkIgYkmbUtIzOwLGABycGxJK6Qsi/hEY4vRZx8zM7thWcS3h0TucM4OF5jNwA3UPi0aEfu+67puNpvP5/Pt+azre1GBPRnSi6wXhbTusZKVwI1Ve7P/c+V3hJpbUDD0cs6/LcM6hpgDh9bO0cpkc/WkAtASCF6gNxb/4HJ3iN1IDsQ7cDkSIrkXEQcj7tdzOvYUE/7c377mv/93dyIxOT1CBID1lv/L7756nys5sdkd31y8/sqj+1zeTE3F/bIlAhvBDFQ8T7w4MJGWRmnPYJWc939oZit8GRE8+AJKYzKx5PZyJ2glJ9q5W+Bi5h3uqcINqdrUa6IK1eyS4Z/gR+NrMwQCRA8FAgA/aiihGIgHDNeuXLuUInb6nw1MTcoDsZRWhiFtVgYT0dJRD+DPq+NnOrhqv/vw+iuP/J//6Y3/7PePiRoQOkytTR2H/Ry83qsu77ILex7XAG93PF0KuTdEKKHAQ5XvrM5+Zh7jMOTXwNI6X1b79YRgWL24q4h59wptGc5Qqe8O1Xcbnh0zv/rrrtif59mvvfZTUy47kHPu+z62LXMgwr7vc72DqovZQghgpqJQubP3AEQCBCX03BsyMyy3jxdszAADs9X+li6/E+onMCiWdAv/q6c5+UdSKTNiTb8xBYMa720hRg6MCP1ikVMPO4Lyzcy6lAgJmnYm+eETp2+/4/7N2fb2NZddth5a66yfr0+nTJj6TlQBMIZuQXMiyiJZck65bRu3RYvKsuaEtL297UHVZqpeiGUKHLxa5mkcCMQUyLPjAcSb8DIrkiJlAwRLKWXDk3k9UL7lF9//U788BnGMGjVq1KhvH40AetSoUaNGveRlZn/xF3/2iU985l3vus7QQiAGMUtsmcEIobRLQ0I1AiQEJkAEImQkZopMTYhECGhMxESBPe+RiEAlm2YC4MAUIoi4ASo2E0AARlMBwxgiECKCgKqqpowZJVMn9MgTp/76c/d+7K++cO8Dj6mBAVpNYbYyId09nThdW7vi8ive/va3v/aaa5944sknnnji+PHjbdtOmqAqzMvADc+QdNzgXaQ89cKRin/jBYAYYgjsTrQQoi8QYiNufK7f8gGAcvZUjeE7v6k6BoNKysqX/tptKefMjGaleZSqItJsNt/YOLV5ZrPrOpWMB0ngPc8BsOTDld3sNTd/X+vatZStmqnxedZf/owVRe8wK65Mex9WW4C2IRE6pdQsxAxoaWePQTfHWuWeXifxUTOAafVQ3eIGd9qjpvvNSTiobnzFy97zhss+es8zFYiaAfz0u68+Ot2vce///djX3v/mK/e/RTOPdgE/MkRDJk8mGTIiVJWY3cbr+E8k53wgYmtmCmrVYetE2m8BNRNnbDVt26MYnIlxsRd7WoKVfmXLewcqnq7cdUcnybIiA0Or8y/qYRcjPCAgERwwUQSGcVmip3fyZzNAoRAQuZiTEWputNVOosudgcpJHzq++f2vv3T/+/A9r7vkt/7rd/7Kh+695+ktAATTysKtxJWs2K7NaoR2hdIru7xyXPX/lmvysk49zOX7rMa0rMjUEEoNxcw8UmYH3/fYm3NkdyzPyB7UGOruGD5/0vRKBQJqEspuBl3/gauv4cr4WbL8UtQ8sEzV+w/2fd80i7VDh2PTEGLXdzllA2MKIbCq+QdjzllNvD2hfyIQEQEBeG3BCGsfWo/p8drnrpKCqUclG3KtG5XCiKkVD7t/FnulyyteULLZCQyIuNZTCaAFAxNTMVNPUbdhdCz6njhQiNn05Ly7474ns2TT9OZXX/ayFqjLhqlh1JT8uaJZ/OiS42bVRccxRm/bm1IGMw4hxijq0SNGhGbWdz0xhRBCiGqaUvLkEKboBwAAaqYASoQhUGxyTkkhS5c1cAi9UUT40M3v/+GbRwY9atSoUaO+TTQC6FGjRo0a9ZLXAw988Qd+4H0pnTbTScsNc0qzgBgCMZYOgwQYGH3uKyEyuWnKEIwACIFDYEImn5JOgRCZkQgI2NRUMGdfDkAhdbC9Be4N5KBpoYu5+1QRcTbbms3ns3kfJ0e7HL7ywGN/8ckv3PbxY0+fOJUK4zGCitIAuQaerq+vv+7669/73vcC4KOPPvrwI4/M5nND7HPWXnNO6+vriNh1XUrJzNq2AXDabczcNE3XdSLi1mUASCn3AMzUNA2aLrpOVBCwUVU1ESnmVSq0fW1tzdcQQjAzqdY2ZweAGIhiCIhIzCGEyWSCCGaSsyBC36dTp05tbW2dPn0m952pgocMfOPtz1asqCvGyV1JGrbHbHTcHbixe18R0Vah0OB9XmKU5TEu8zdqDWBPrU7YF3FiY1ocvqCaPenAWYWALBmZmZcfis9TzTlpNU2jETmKBVAc0of3p60uH2r3+y+H/+T7Xvvxe57cTmWq+ysvXP/xt75in++9/5nNDx178v037ttDu5RZgcPL5GIcSjGFZ8ngNId9eUKXagJdeGgChQ47fyRTAGLHssShInfnyxqY2kDrk/iy9ebpU9sPn5wDgKnzJUB3VKsiImrl0QAlSQCrjdrMTEwLmy3rL+RMoRBUA1M64N1kZmBashh8kJQzNRRu1ByeqSwt/LWcUypO3icVSodAYr7nidMH2g0AuO7yw7/xX73jMw+c/IPPP/bp+0+U8JgSG1wotzpvrj5kVa0JIvVwzlopVmBZWP/y9UqzKwjeVQgrp6LOTii9IVczglZ4/eooYubKqYdht8coG3j6WQx6x6IVxw5XG6yEQBu8wNA9++Gyu04GsL/b33x0GCCo5WxqKmAxxhhCvUyKiCKQUkZEZkopiZoh1dB/bZqmiREAskhKCZFCCJO29cimlLOZEWLTNP6xIrVbQOnIV5+KWcRUAZGZkb3QWo6vgGYvm0KB3ybDmTAOoZ2seb+BvkPVbMssDhADVYU+ARgiKeh9T5xadBkpvPE1l199xdWNdlF74FC91eUxTu7jrqdXFA0IiQEBQwDmEEoN2GcpGVHOqUupl6xqfnIQKWUxqTE0SIYoAijCIn3qswIoMDGIMlA7NbQxDHrUqFGjRn37aATQo0aNGjXqpa2PfvSWk88df+CB31XQ0DYhkuQFaEKONbyAPTwCCWvkMlqZbu4WUQNANEMzUCwkyL9tI4LnbwAQqIpJ15tm1BRSL5LFRAFBBSWLSEq5TwkJzSjGtZMb2w8+dvIvPnnX5+7+2kOPPZ0rMnCLHgJ6ILMZxNisr6+//obXv+Y1r0kpPfvsiWePHz+1sSG19Z+IlBBMxMWiSympakoJEExLR8Gc82KxUNW2bR1K5iyIGAKn0mlQnF32SaplrDAmInKm3Hedh0pjdRRnkb7rEDHEiABaU6crCCiAarHoZrPZcydPbp45k1Jf/IcGBvoNCIFY1Tm6Au7vrfvRC9Hn4Q+VQVdnJq26v3dta8cqEACQuRgYsbj8qPqYSzRH7dYGpgbew3IFfSHi0N3Lqm/7QOf+ls888lPvfNU+GfSlRyb/6G+99tdvu8/3/2ff87qw73SI//u2r+6RV/u8shpW478A7AiLWP6zmp8BoNhXD0Jsv/f6y773+ssOtGOr+rVb733o+BYUm7ADTVnZB1WxSjoBET2PAsxbeO6Vj75i4rXqxj6g3DiPSABqK+fKln59VSu0d5lpgYhiCgAqfgjLEBkFu/PB40k08sHmNyDAu1570btee9HGvP/sgyc/99DJux567vGTs3JY/jRERB/wg6N59WDOdZBQSwIAxTRNUBi6mpnhrnf6siJ5+evOoVKh8Nk8V1VW0jwGQ/uOPURceWXFOb77GJapPDs2c1bd7uy9t9VN7rXAivB5/zpsulJ8AdNkpipZ27ZpmkBBVbyFpZ8u1eJu1uruJ+I6jtz3XTKF+r4XKWkVAKAAKWe/uGVGg4/9Ff+742wESjmDgHcmLCO1msrL0AUAsxJyUU4KIiYOsZ1MRNSy42kc/OOlJwSCARrxmUV+5PjmZ+97kprJRRdfura+digqSw+qUGpIZmZZBQGJOYsnZ/gnJgHCcsDVYBBVzTmV4kodPrWvI6iIemmKCImtlKVUpBXRrEDtoSzSq/WSj/CZLGFk0KNGjRo16ttDI4AeNWrUqFEvYd166wdE5czpk71R04QYoO+3TDIX4x4oewQjAoGIZlWCEu5MYAgKIoxABEGI0MgMwAhLEyg0QzUk5MAhBMlpsdiWnJh0raFue94ttlPOTdvGtlksus2t2enNzUsuu/zwkQumzaGvPHbfZ+786kduv+vp4xuKIAbm7Q1rnGdxviEcOnTola94xXd+53dOJpM77rjjxMnn5tuLtm3922x1CmrfJwAAMBVVs5STmSHgdDpV1fl8vlgssIZB55wNwA3Ls9lW3/cA0DQNczDrsH5jLkuaEXMTo7cTNDNm9iAOEen6HgCiA2jVlFKfEjP1fe8ziVX1xImTp049N9vaKhAACcBsmf583pD4+bVCIr5xwl0/7KmdB4oIFF44LcEvhCNmwuCGU7fSI5GZKUgxAJYk6JJS7H0mHa4BuO8ZzUqGAAGB6UFPzamt7l9//P6f+6Hr97n833/X1R+88/EnTs3f+uqLvvu6/QYyfPr+E3c8/ByaHtAabytGSI8iofprBdLFO7oCnYuR+Zskz3v23fDeg0tg7MWeoWukx1VbBa1abM5QfaAVtK0clQ5M6yAyMPEGq1io5ZAK4kEu3kzN8Z1Wz3UNswYoRNG9/aZlV2fb/d0PP/f21158fifqZWvND73xih964xUAsLmd7n9m85ETW4+cmD1yfOvB45tPPjeXVTPzqp5vQFd4jmiApFRf2HsuQsGgJoW3EwMuE5mX6zxri6bFU1vg+K64DEQsCcX7KX7Y8glZTjjuRsa1sLTnG8tvsHtf/KWzIf5ePNqGBHLw6y29ggESTyfTtmlVRdVEFKoNuWkaQMxSbr7V3KfAoW3YzEQkpV7NEDDG6KfFE6VLj4GytmXoMwBwKX9QVlEzKWkqWCM4qHjyDRGAiUIMpiaq4JXalNbWp+100ve9qqgKWEn+KFk6JeIFkUgAznTp8195MjTTV77iqguPXr52wVoLiSSBZlNBACTwvgshNF3q/SNyMpm0kwkipJy7vgcDIgoh5Jz88zTGJoRgpkhERCklVWNiESntHJmJGYglS991pfStqhhE4fR8dnpuW93hQ+3m1qnpLT/5kz/1e7/3QmNp1KhRo0aN+pbWCKBHjRo1atRLVbff/tsp96BN0txOmkmMAD1qBCBCJGZANAMRU5WcgQCp+leJOEtvOWPO2SQQxLWJmfa5JxAC5TK/HtBwMp20HFUl96nr+qYJMTYUMc8XGcPkyJF2OuUYE25N41p7wWVHLrxk0cP9Dz556yeOfeRjd5w4M0sr1joDIOTqDjYO4dJLL7nxxhvf9va3nzx54oEHHnrmmWcBcNK0YBY4hIYrsnLjlCGiB2j0fUfEMTZM5LOemTkEJiJRySoiggAhBg/ZAPepIYoIlKZc6DY0D3HoUzJP6iTqUz+bz5omOqUiQkQTySlnZwpkIJLNtOu6zc3NM2dOL7YXg+UQYJj4/PXQYQTb9faznbMIO1Niy3new6FMe+zL2cbIPTaHANU7v1yqApu6NSrd5crv5pRU3HoPlYL5VVBRpMEfXagNAhKhamn9hoPvj7ka1aGAZiRUD1WwARTWSIriXiX0K7z7dD2vED7w+cff/+arrr388H4Wj0w//97r/+ff/fzP/dDr9rmFLPavbr1HcrKD0Wd37+oy8MAATAZEWvbep9ZjtZyCmyO/UUHYe8hMJTkzHmbxD2kQ1alp4P7H+jIiAjEi+oSGEoKxhOoAYCW0/sBnrZA7d5riilPcN+f7VqpcNXd5xU1cuF/ZZyhlECACsA/f/dh5A+hVHZ7Gm66+8KarLxxe6bM+cmJ231Nn7n3q9Jce27jvqdNW7doVTpY+qyV+AYGo9hIUBQRirqUKN5tXO/RqnLQaIjA1HiLh/Tz1LFiLAIT1ghqYldCe3f0Jz74wQ45I/bvt/gl2lBPqzIkV9I7D5Tp7G4Y70sD92qnt3g/bBZzPYurVrb+zzkakaml7sWWYp7K2tjaZRERcLBZeGmFmROKwfP54tRRLfwL0j6HQMyAScQzBzLJkEUUEprLziKgqABBCrAXXEsQCCFoyptRDOUov3FI3FSrtgr0JITjbNTMOTEhHX/ay2Ww2n88kdaZqamhoq6EtHtVhIABfeeTpWz70qZNvv+bG11x6+dEp5wXJIqBN23YyaUUSEsWQRNQHYEpZZC6iUpof+J3UQ7llUdRKPFYWAPBJSF419M4KKgJZSvNeqCeNGQwghrW2TamfCZ5ZtN2Th+iCDkaNGjVq1KiXuEYAPWrUqFGjXpK65ZZbZtuyPt3eToyBY4iApmqATExc5raDU0ADRQBwFFj9hJ57yYgBOTIylAZ7kYERyTkHECLHyIFQ1Jipadt2EmNgJovTNWgn08NHQghgENeRgShOZj3c/+iTt/3lnX91x71fe/ipwYFpxR1HNWhVp9PpRRdf/OY3v/maa65ZX19/6KGHNjY2iDjGyMwi0sSmaRqpk3a90VwBJaLb2+zRzwrGkgHMgzSaJhITEolIjLGJDRho2/q3dzPo+4RITGWWtKgG5mE+tZ9hb/sUQqg0AYmYA6upKgVEM0ip397ens9mm5ubi26Rcy6JzwfHZOfWC/PTOiP7hZfb5abcC03uJra7AjeWv1cu5HhQB+ruJxKLqxR2kqaB9eFKOKyZRx0U6mdDpi1C8e5Vd2JtY7fDAukT4RFqMjLucRwvLLMs+Vc+9OVf/+l30v7e/93XXfq//viN11x2ZJ9b+OCdjz74zJkKYw/mgB64su3I3Biuqt+zq+G5Oxf7xouxXAgovFlrqWIHOq64CocBMJQKlrZjWKHPhUGuAMmDCVcGIA6e2J3D2ur588pGfd/K7pSRWVspfvRLT/zs+264YL09+P68gJpA115++NrLD/+dm64CgM1FOvboxmceOPHn9z5zcrOrRB+XIQcIyMU/q/UoHaYjl1Lf4JJfnhQ09McpIiASEwAi7Tq9VEpNOKBcA0PD1RpXdSjjyrVerYq5L37Y8HIf6pnew+K8XKRertUFcMevWK7qHnlHZ/Hn3VEkK4MDdyxoJiLdYmEGROWzpmma5UhGJMPBuawKAFpOMyEiBg7YlrFORKpKShS9nSANx6FKAKV3LgCAh6dQKcINALqWHshzlp3llsKbmRkECr4Gp7whBgUwhG4OOSUVsbOTUQwABBDBjp+ezba21yKkbvum615+OMgEcoOiKil3YIpIRAsE8sBsJALAwVlfwb85lwcApB5weSd5n97ylMbSmwIB+i6ZGhMTEzITkQJIymC21jQpJVGMr93UOX3gf/yhv/crH9lziIwaNWrUqFEvCY0AetSoUaNGvSTVtjjfYgyHiUPTRIVkOYMpucuZsHzPtvI1nYb/IjD6D8QhNBjWJ00TuE+diiKHSRsCI4MBMXCA0GDOkHIIvN7EdSZgBFAUOTKZQAjQtLnr82IxXTti3Cg1X/jafR/52Gd/59//yXPPbeaz9hsRkd0sJioXXnThm970pve9731bm1uf/9zn5/P5pJ0cPXI05ZRzVlH/wt/1nfeaU1MErHOXYTqdElGIIUn2b8KOL4lQ1NS0zllGkSkRtW3jQdWpz6sJGymlyWRCzJKz82gRYfZOU2W69AAdYgw5R0RaLBabm5vPPvvs1tYZEwEkADSVc2CUl7B2m7D3I58x7hAHAKia0G0nNS5WdDMREclExMRApKoqYgCEREwiGQyQSEXd5uv1EhussiubgCWlNDiI/1dFct8fe+jZP7nzsR996yv3+a73vnm/vQS3Fuk3bru3phwcdKBY8RS7cMX3bks+6rRx8Keb6XmkJp+3AjMCIiAhK+qyGGNa/bdYCiFDMMISaZZbeFlQGYJtl9UTg3N3tjynhlqF98cEgpUkDyvuZhxszsVtvIz+cJdxgXeDmzsl/bd/ef/Pv/8NX8cJ25cOT+K7r7vk3ddd8gvvu/7uR0/98Z2P33bPM2Xexq7YcSQyNUmZ2NP/y1SDXGOIBxEv6wBUDelnzaUwb9GoamX6QnWLn4WYhzpDKRetTHk5q/Bw1t4i1hkSy/6HK0WpspXd9Bxsr0pZ/djbvcXzrglqzp3O+5xU9fDhQ96f1p9XWu+tCqAt5zIRJzbRz3wMwQxUtU+9tx0MIeAQUbKyqymnGigE4LjfAACImZGMUEw9wYNDQEQOgZkQULOk3IuIp16snq7p2jS2cYtpe2veLRZetcNdEN6fkp3o3V95HLJedcWlaxcfmq4dCnmRuq3Z7EyMgQA1K1Eww5QFmTgEql2OU85qg/sbVC2LiAoReX4XIqlK3/eL7W0RadvJpG1jiKbm/wXCUk42EDMFyKKkWZIpAjZZCf7gl977E//81vO7jqNGjRo1atTfuEYAPWrUqFGjXnr64J/fAj0cnRCGyG3DYKICaETISIGJS8SzoZnzQzJrmJsQuHhEjYki8TRQRCTUlhGaBkMTAhEaSi5f56UHFUAFZiQFkNxnU0EzDqwZujMnwZAoYOTjJ05+7eGn/vjPPv2JT33h1MYs5V2oyMBAzWD90PpVr3j5TTe95brrrnvi8SeefubpjY0Nn07cpd7MkCgwI1FWEZ9WDORW65SSNycsk5RVmRkRcxbm4CyAeMhjMFPlwERkiN5NLMZgBp7FiYhN0/g3e/AgTiJEDIFjZPfBuePMOUwIERFPnz6zcerUqVPPbc+3VRy3DK7KA6fUVu0RkLG/xfZaZI+kjr2W24sIwb55DVbwuVw/Lre1+1yoqLonX7T2XavuxcIEUc2gMmsnkCLZr3ahNmZItgTj9SDcQ+2vFYYIcH749f+69Z7vuf7yl6035/He59H/98kHTs97Nwge1KJdzK71yiAgDD0XoRywVYtjIanfdBEVngje8ZRwSXd9bGHNjvBwb6p29noM9fAK6R0c0LUJ4IGvZnEJI6xkPMPKCqHYxodAjvrCEtPhckxXM3A5mj/4zCM/9vZXveriQ+dxrs5DhPiWV134lldd+LPv6X7/s4/93uceW6SSXj1MCCiTXIiwHDJILc4t4SYAIFp9FZYIVXcHa6j5TYWSMkBxMg9gd+WHsmYEBBrM97b6iNkjEsdMPVgZdlhzX/hcnOWHtuGVnXQVrbzi3vl67XYY6ffcmg1VIjMzSzafbanq+vqa1yNzzjV/PvhHFSEwkXKZWOO00zeWAAAgAElEQVRA1gC0JGOU06WqIjIYkCv0RzNdsVZjeTwCmogBmFrWDIBMpFn8sakZzUxyRkTmMFT7wBFwzrGJRBSbVqcKAKnvVbKVVBJcrS0agADMRR98+tSfffzYd73p6hteeeHEOkszkMXUmkCMtuwMmVNOOTWxsQyqqmCIGEKYz2eePR1iE2PMZnmec85t0xCzmrmXXEXms5mZpT6DARENHxzEgTgAYRLpsywWkijEplD3/3jzj/34zX/4wsNj1KhRo0aN+tbTCKBHjRo1atRLTLff/h87kdSoGDcxBkKRHsGYMDAF4sAUCHEJoAHByKwNPAmBwExEJUemJlAbGVVMhFGREAMbgah6OCSaYe3kZiKaRUVUMgAQoCTIOc02zzTtNE4Pnd5c3HPfYx/7q2O3f+yOe7/2uMIQN7mUB08ePnz4qpe//DtuvOnqq6+OMX75S19+9vizi8WinUyIuXQoImqaJuXsLY8IMXLwLI6u65hK0DMiMjMFFtG+7z27w/k1YMnEBERmQkHpFjllVWtCoyLFmcscQ0g5m/n04QJiAMxtah7KqepR2hkAcs4bG6eee+7kmdOnz748Zx/xQbUfargfTo37W9XZ713lSgfyDO6Yu45oxeG3wyZptUmXA333s7v31Rcg4mLdNfNp6qigZqZKfmm0Wvodnex0VA4YbmCMtJK8cCCd2e7/n4/e+0s/duN5vPdceub09n/41APVKboH+38BqQ3QCgqs9Z8quyuYrULbFRPxN01ENYKj5HqXsoxHF1vJEl+JH1EbqhRDvog6vvaqBpYs6ULdz8fK6v5O3w1drmcYGrZSDqi7VV4v/xuCCyqUNPLh3Gf7337vzt/6mXcHpvM5X+eriw61//gHrvmJt7/iN29/4E+PPQkGq4nbBd0bgJkMudc7TtyyaGOmHotkpch2tjvWTEv7AC/veOLEwONXbOww/DiA1D0ehzs/EfbY4vloOYxWCmB1Y6tmaaujaOXNez60d+TbGJh2i4XHN8foft4C6xVBwMjIj8XTxrVXM0NCNfOJNVDyM2qkRsXNHqkB5UPHg+trE89hLoCBmpeZ0Zj9jHkiuq8thBBCGHYJCUW16/rWtIkNIIYQrTUzy2Aq2VYOuhYOTAE6g2dOz2Zfmq031JBccbRZjzjhhkMTQ2AgAFTzj/+sqkgEJWS8TEChmk7OhDEEP1CFjICMxIwxNkTUd11OWerUJQR3zYuIhAgBCQxMxEQpUDQiCqiGk0YWdssv/ORP/erYkHDUqFGjRr30NALoUaNGjRr1UtKtt96ac9cG0B5iwwiqIogamQJjZIohMCIjUEkrNQBAAwKNiIyGqiJJUwcQkdgEVEUl5dxjD9SBkIlITp2JkFkkijEwUZ+6rlt0/WJtfb1pGkCezWbb81lK/RrFDvrP3HnPbR//wp/ddvepzTkzMrGIquwggG5zvfbaa7/jO2664Q1v+OIXv3js2DH1L9Gii773r69d1wHA4cOHu66bzWaIOGna9bW1rdlWTjnE0DYtIm5ubTJxO2kNLOW8WHRt28YYAACJ1Gw2mzHzZDoNgVNKs9nMDJh42k7AijHQg6HF0x6cnwEAADMxk0+4FslmICLb29uLxfZ8Pt86c6bv+5Vv8bSc5v83Yj39urV7dvzXK4OSgsIFSaioM5imCaJum4PSXwuQiDiQqRnY0J8QwEl0AdOexO3YZTWCwsFhQW71quBBMLwLK1pDxD+567Efeesr3/SKC16s8/HrH72372XYwwNXKnayOqzZFqsJBw7hrPqNh/d9vbu+b5GZSkbwbmc1CajQZk/RGfikDWyv2pSXdF2rNR6B1KScs9L+7oARHAYV9vm4sOLCBgAHdhXarrxFq5MYAEBr7PiStrpnHwwA73n0xC//4d3/7O+95UW/gV5QFx9uf+lHb/iBGy793//gCye2UilBEGHNF7YaYgK7RluxcpuBZCBCZlPdGdVcF6tIsXQVrDMkSt7LzrgM2DnvYbXKsuLAXu7Oizg2X2hNA3Pf9xoRvJupPxLMQHLa3DjFsYlN27at02QvkZpZzpJFPT5IsnBgZsopiXrdVoiQmN2nLFmg2p+9iaBkRQRm9g6qXsjxUYqASB7VDYPNmZlV1MxCDCmnIYTKtLRJkCxgpilnt0jH0ECLCN1ClvMpVk6NgSVn4gpfeuBxy4vvf+cbL7rk4ksON5MADWFA6rouZwEP2gBIOSMgEqackbBpmosvvgQRu67z3qeIFGNsmkYki5ohiGQVgUOHykQJD3nxW9RDPDgAkoiIT37iRjn0i8Wp+bxfLLQ7nOTUb/zMW//xb96x7ws5atSoUaNGfUtoBNCjRo0aNeolIzM7duzOZ5450fez2HDThiwZQQJCRAtmrApJDUHBRBVNibCkcKgoQAbIfQ+qiECmoNR3RoXjIRNhoNx3ScQMmnbSMJOaSs59UjWOzfp00kynCJi2OzXidn1y9JLnzswf+OrDH/7Ysc/c+bUnTp5WJzRaqBEjIyECZJGjR45e+fKXv+Wtb73qyqu+dv/XHn/i8e3FdowRfG6yuDXM1AwBu0XXp2QGRKRmi26RUlLVACFLLm5q05RSn5P7l93+vFgskNwkTQCQ+l6EwMBDnxFoQCHMrKpd33sEqqoOARQ5Z1XMOTtiQISu6zc2Ti0WXUp96jvVsyYxP7/Ox9qMexHUF/JYn2VNxJWXd+1DdXbuSZ+xtjGDXeZOIhp2ZAiORQMKJdQVERVLx0gi9NjYwkUJHTf72ERERSTPDiUSEJ+RvZyQjlAbdlVu6eCsnPwhvQEG4HbeMjNTgWom/hd/dNe/+aff96KYW+95/NSH73pk+BXdJ34QBn32oqshxmWV3hsOlk0a/fVvJoBG57VmBog6xDxbpe4VBMNgii4HsJKHa4NnF8E7g9ZD0OWfDyDTZWx0XfXQ5bI48K3cyMtdKyez7P7q2+seD79+8PMPHZmGn3v/m7/5DBoA3nXNxb/zT7/rf/oPd9375IYHNhvaairOwKBXZZX8w3IhWNLn4eWdIco1E8XqSVk6x1fOzcqbaubJHtdsuUt7XtBVF/My47yu1fbIsBn+es4BMoDWs2Z4ICCdY1wNER7gw1jUDHo1VUmTdjJdW2MORKgGZbIOc/nIICqp9IhmllImJGYyAJ9/U5M3rNwZ6viVygMUoFTpVAulJgIwVROfn0TkY5iIDMBMh5KATzHJlGMIHl2BRN5DuG+ioklKKtmH8HB9EKBgZbNnN/v45MaRrz6GgQ8dvhJMQbXsbEXmfqGJKPhWCJm5bRt3QmfJXllkJr9WNaTFU8lLC80Qimk65yyq6G2UibGJbskXJKAmhZC0n2Xp+fSp2anrH5sZ7P48GzVq1KhRo76lNQLoUaNGjRr1ktEDD3zlxhvf8pGP/CEAxBDNBKwnAkYIBqyKomYmYAomKYFZYCIwMFXJjEhg3faCiaaTiX9HziIhhBBjCC23IQQCETBjDmuHD01i1D4t5lt9zhyaydpkcmjNmPtFl2cdtWttaOPakccfuuf2T335L/763oceP67FZQioBmZUZuYSEsWmufKqK9/5zndd97rXdV1311139X1/9OhR98aKChIpmIi03CKgmTGH6TTEGMFMch9DRMTYRFVV08lkAsUYqsy8vn4oxiAi29sLBGDmdjIxP05ACtRO2mLZU2dQSEQe0xFDYGatKRwioipmDgok56wq8/l8Y2PDUzgAzsU79vxSvC8n7l6ZDHu98fm8yjXBGRAqNl7CoD3WdM5v8ZUqF1Z61lJEBIim5mmz7M5xNfbp+QA1rACYCAlNBRCJnZiAqDplMQQAAsRQ36gFYDlMtkIBCUqGQIkJKODEsF5LsyUI20HPznmm9papqtTkELjv8ed+71MP/IN3X3vAteyhX/2Tu9XjWasQ8dyk7Bx7t9NBitUFXa559VUPnN7Mc6IP3rXvfEXLCOrVvS3s0q/hDlfs8I+lBnZpy5925CYc7KwZgJ3VtxCHQOnCVK3i7+rK3Lkh23HPDS7hOugMAP/9J+7fmKVf/PGbmvBNzeJwXXpk8uv/6B3/w+/eeezh51QygNV2i2X/zyGvEHKJ7EBe8vbVG8fjIJZrwWWlZ69q2I7nk2eDABSSu2O1dYis1B52bGL3rg4zB0wBl0bv1YXOPuCzd28ZFr2LQa/u9iqVHezc/sEGqqK95L4jxCNHjjZNEwIDYhbxTyJPeVYzdBbLDIA5lw6rVmOdfOXL3IwaP45I/h/vdgBDkY8KX/YoKqjPkOHtQ1Y5IppqSomJmFnKpx2GJsbUGNpiPk8L8KAtWLnXfNAktc0eHntuoV9+pGnbCy44evF6OBRgAoKa0fNOvL1pnYXhEUmq1veJqFjCDcxUck5dp376dDil5UNWA4SAgZiyioggoKkyaYyREBTQVES2AexQExe4SGAXHb3we37zji/+rVfDJx6CUaNGjRo16qWjEUCPGjVq1KiXhm677QOnTh3/yEfuMxNkVuml7whVxNOKUcEYBoqphMDedbB0o5KGuQlsRyUQN03DBAigYBQixYhNIM2Y+8NHjhgjBAoGIEIE7WQS2wZjpBggkPRJkmBop0cvnPVw7NhXPvSRT3/4ts88c+J0YRKFEigAqE83VolN87prr/uOm256xzve+YUvHHv44Yen0+nhw4eZ2Y1jItK0LRKJZLDKGqrBSkVSt/DUYETMOZtZbKKI9ClNptMQQ9u2/t2+aVrvZ8ghgENF05xz13XMHDgEjowEiH3fg9n6+rrPd/Zv0S5VZ9CWc+77/sSJE1tbM9XnYXkvuh9rX9j6mymsNrbqU1dEJDUIAGoqYkOIdjWzGxMRpZQQwZhNC0ZexmcgIEBSAQCwgmNU1Aqjqdtd5k2s2JxNbJWFwQ43MPr/DmKY1WVMQPn/X7/1S3/7zS+/5Mj06zht8LEvP3H3wyeWBBaHDRzEAb0zSAGX/1fiEOpPg2UTKyr85jmgmXCFiS9V8TFiZYurJQPvTTe8w4a9LztvuMLIzisrZhgWULk8rKRwV2/+ig+4vmFpi3a6tzzXDmZh4On2p3c+/LWnTv0f/+CdV19y+OB7+PVqreFf/fs3/czvfP7BZzcRkUPwYo/tHAE7cihs16iqCw3yJyoQIQX/1dSw9npdWW6l918diqaGwxvVVHWVig9Vij32YPeAHVi6HxHRWdeiLOUTfnDVXr2HbIhc2fFg2bGi53n7oK7rT558rm2bpmlCCEgIiCJSH0BoYKKSRfxJpqQCIqUnobkJOoQwzL+BZQxNSdsYfOYEZGq7i5Qevjxw53pU4F18mRgRkwgwcgzI1LTNocPrZzZOb22cnm1uqu6oipmZAiiAAGi2J051d9z7sKTt73n7m1558RHUjtRAsmkiryyaiUhKSc1EvV6bzRSRmybGyP5JjYhN0yCSx3e4HdvURCV3YottVc0pI9Bk0mYFFdUsOeeck19xI1gIzLq+F+LAv/tLP3jZo6f/3Q9e/1/c/OH9XKlRo0aNGjXqW0EjgB41atSoUS8B/dEf/VFKevr0CTMNbSQAywvURAxoYgCCCEgldRUAkZGJA4cQmYkJwDQgMmET2hg4UkBTQDUEZAZS6WfSLbTrwrTByKbYL3pLic0IkZlNRZNKBs1iihQnG2e2H3j02Vv//NN//dkvP/TY8bRqBV6Z/K1mR44cufyKK974pjddcsklDz/00BNPPHH69OnDhw6HGJz2Bg6AQGU2buP+YzULzCEEAzAixqVZrGkaT+tV1RgjBQciJiJENJ02aiqqgEiIFCMAeA4mAAbmJrZgIDk7dG7a1tN1B/oMZkRoRn3f932/ubm5tbW12N4+OMs76ERh3PXz3wyD3nmkpb2XDY7p6kUGBCVFJffDKWppqFXNcaqmJgBgBiqe8+nEp/giK3scMNTAzIqFbsjbXYKqlRyHpX2y/qW6pwFWGiGet+Z9/tU/OfbP/7N3nfcakuivfegLsLqXw44fTOd4x/LAq530oM7qF09MuLcttmiP2+F5fbp7vHY+F3SH2XxfNxTucb2G47Lh78tSAgAA3Pfkqf/81277h9/7un/4vddNm2/2t4z1NvzyT7z5p3/7s4te/Y4qybqDhbfcwkUDrFyN3wYA3Mk5C5Rf3nCGe4DQlZkgZ8HkuuaabuR7stwJ3PnCjlWtrKXusdtvde9Mod0MevdgLG/EA9+KtsMPDYAqebE9l5xS34UYQ4wcQggRvJQFPskGs6iqOgsGgAFA+96KZFUaop+WTL7sLJJHb5eLiY59oR4kLN9YPh/NjAgZiZg9XVlMQElFGAEDE3MIMcRIxEa2Oj/AalnMAHq1M508/MymqBw6cnQ+v/jKww32M0gdqIQQYuDyLv9ohjKjCMCYg6n0naWcPC1E8oQ5iC6f11kkp+yR9YiQsxBQSj0CmVjfLVKfRISZAE1AOmM1CkBg3Ag/dc0lU8EP3vwjP3LzB/d1+UaNGjVq1Ki/aY0AetSoUaNGfavr1ltvFen7HhANGGMIoJ2pAmIAcQpiSIJsREDoGZIUmEKgGJmQCNDUckoqLTdMRKBgYqbEYJK16/qN57r5THKaHppS4KzazReatZ20TWw4REVQBEHg0CJPKLYPfOWrt//lHX/4wdsff3ojZVAslsABnA5GwSuuvPJtb3vbjTfe+PRTT//+7//+JZdccvTo0RBCcbyqMXOIoU9JTJsmqnujckbEANB1HQI0gYfv7dPpNDZxPp8TUvv/s/euwZIc15nYeWRWdd97B28QHBIAHyIgigApkpJIhWRppVhqJTGk8K6tpTbC4QivN+wNOyzZUtihX45AbNjhXcm2vKsN21qtYtdrrb1BPSmJIiGQBMUnSEMgSAIg8SAGJAiAGGAGM/fR3VWZ5xz/OFnV1X17Zu4MZkD8qI/EvX2rqzOzqrKyp77zne/UdayqlPNsNjMzZo4xtDlLzpIzM7s8jZk5cM4ZDAKHtmmapjEr9e44BFNtU4ohuDLaxXqz2ezUqVPf+c53UtuK5CMq4zpYV47riJ86LHneKIJ+hehF6/LQD/NBRQpddsChzrL/FAAws6ho1lhFMOjdSzz53VXnxY23U8USlsR6HZjYYnGLHlrBFmHgYU6z+0whYi+V/u9lrvaxr3z73/+h5997200X09ISf3DfN759ah+6M9PPoEsX8sKSY+6mV089w/AFXKJe+NJRuLJNHHRHIa7Qkf5O/wM2Tbc1hvISCOiNXOVSOz8Ilx2S0Q9lvdaPEld+rYjZm5R+52MP/ckXn/z7P/nWn/vBN269sjT0rddv/ec//uZ/+pePZVXtC336YA+JhTv3f7CuENzGPT1WpL1gWVWdpF7ZaQON66pezxpxv6O+l43T8jxz1Z3ZO+W1gRoQAm3efwMHvfo+rA0WAQEvOK868nlIXKtaSiqSCANX9aSeTIjYANqUVM3Td7yQgIUVjhgAYoxImLMASH/4a8MgJCYiQDCQLIBIRiDuIWXghYbRzExEiwRZlJlDYFfBq5qBKYAR1nUtmRrTnBMRcYimKgMCeuiVbgAJ4MWZHDxzIPrQqRdufM/tt+Bij9KcQOoqVDF4pQUkNIBYVVtbWzFGZg4hpGaxWMxTSq6ANtEQI1JwXXOb82KxaNuWiGKM9aTOWVQVDqAKNRMvZnPNGQx4WgFaTi0QxzjdCnVGVKNjC6AJJ4UP3vV3P3DX75//2o0YMWLEiBGvBowE9IgRI0aMeFXj3nvvTblhqIgWUGHgmNumbfYZNaCIKBFSCCFUxMxEgYkJmTAQBsZIgGhoYCqEGJjBrG3b+WIhqTUTYkipkbYhSQGxriapTZYSIkZmruqqrjlEZDZEA1RE2to5vdc88dg3PvzRz9/7qQdeOD1LWh5c3Tt0oAyErcn01lvf8O53v/uOO+74+te//txz33nt8deGEFJKTdv4szwSsnKWnHJSg7Zt2jaLKCG2TXNWJIvEwNNJLSUtNzdtE0JoFg0gcgjMnCUvFgtVJX/MdusPkc7Eg0VkNpsREVMIFHpSomma3b09L5PkfLTzJk2zmM9n+/v7s9kste2age+rGQZHroy48eOHGaLB68IvEgEAECFC4bEQiKl3jkZCBAyBSFHZQgjgNMRydnBRNVvPD5oT0P6KAEzBUME2kIc2GGo55tW3cH370Y59VQrab/wnf/zAv/vVv1V1ir+jY3fW/ot7HuqatBXd5UWObk2Q6wMbEqaDVx2VOsjiPyK+8Pjzv/OxR1bJ2AEBvNqSCy1joCrQziQem1ZPv7hfRrCuF+4GuHTeWBuVDV6sdr1GUF8slidgyCav9bih9TUh7+ofh6/GCl7Ynf36h770f97z8N/+oTf9zLtuvf34NRc97EvFf/iDt/zJA89888UDJCRkRCueQmYrB+r/6/IQiGklBjAAIffhJSQi5k6BC0sfk6UkGrF4bJsZIGHgUBp1450u5aFcW/XkkwuAY3Qu1b/v4mSSs6RBQGvThxCKpQQMpk+33Aw/cYkRvbLSqImKYtcRAhhSyjmLqLpfCCJRFnEzKCYGADVrU9sP1VQ1Z7O+uKKvqZ6OA9R7QEPnAe2VCRER0Ki7EN285sAe5PMgBIWAoCLSLhYtAKj4ujCpq4WKlNPoBHtZn/s7xBCS2bOn253J/nU7L73ze99w641XR0jBhEBcbU2MqubVBUOIzEyIZjuqHgYx6OrWljAGAgKIimQR1RC4qidtanNKkiVwDBToRgQDUBUT0ZQ1VdOtECdqQRTOHuzvN21uF7m6Zl+md91111133XVpV3HEiBEjRox4xTAS0CNGjBgx4tWL++//7f3ZqQjXz9NuqDlWQdo25RYRQsCIzEieTxvqmogYkQmZgMFAE6iqFD5PVQKRMaUmg2Rtk6oAqJhlAcMYJpNYhRiobWZqQoE9nZhjXCqzkJDC7iw9ceLZj917/2c+/9WHH/1WdhLDC1UtuUdQs+2t7Ztec9Mdb7vjxhtfs7e39/jjT5w5c+a6665PbZrneTF09hJ2ThV0Ism2bVW0qqq2TU3bIGIMIedkqq7zSpKJSHIuFphUHraziJnOFwsiAm9W1Z/Vs+SmaUIIgQIRE6DnR4toSqmz0CziXMl5f39/d2+3WSxyziVJeaO1gF0yk7FOmmyW655r0znEf1a0iZsqGh5hDLDKNrt1wUBAeli+iwDorA4ONctLmWHhEP3aut7caUjsKKKl1Wm3yYsRdgXtOpvYYgANsPIf9PYKq5pnK8YdRzkNPVZaWh7306f2/++/evQf/M23XVRjAPC7n3hkb57KKYF+fCsk+cUObm3T5VU4nzloHnzqxc0E9Bq7vcS5hrB2wwwI5Q2f2Li1P12b+O+jAjfdupdIOl4MbHfW/pu/evTf/NXX33zT1T/+fcd/8Hte84433LBVX9mnj0D4H/3wrf/Dhx4BKLcuQhdeGxy0k8hLZ4uVen4rym8EcuEz+tLuRRtdIkse5Fjeg4AlA6Kb4ogds9mZUuDAffsCGNhtE6CBCiAyc6wqwJSXQcFDIufi6uO/hrpeGPCrK4eMeAER9GooptvYmWZ0NkFmgCFGZ5kFRLISeR3CYi7ua6CJWHdoiGgAbsxRYnsAZsCE4JFUQELkwODfaOJWFuXseIwOCYmIiIkQDFTNJHstRDI1AO1Npk0JgAD93w4SQqm82i28yyUfwcCy2ZlZfvqF2VZ16uZb33jL9JqrtznognKD6IFpM1VVE7HAgZgQEKmiUiWyLMymJqIKgIghduUZ1JCQQkgpSc6mSkCEHLx8BUCTmiytgVTTKXOVswqGGEnPvNQ2SovdRyZ3vDZ96zwXbsSIESNGjHiVYCSgR4wYMWLEqxRm9sjXPwXw9RfOIMcqTirTnHVRTXi7uiqQRYJA4B6RxBHB0JRMSAVNFge7khsufgagalUMFuMiS2Cqq3p7e5uIk+RY16GeYD1BUJAU0wxMMBC4L6UqaLacZL5AZsPqicef+NjHv/iv/u3dL+3OBAAQCLAzUkAAZA6AYDkff+3xO9525/e/811PPXXiox+9ez6fMbMZtG0rIsQUYgwcVDW1bUqprmtmBoBF04hKXU9yzpJzPalTTotmDgbEVFV10zYiEkIQ1SyChCGEuqrRNCedLeaBQ1VVVV2rVxFMLSJOJhN/VA+B26Zp2zbGGEKoJ9XQl1M07+7t7u/tzQ4OnPjseZABQ0GHrljZZfBiyOMcpjw28CCH+A879DlEZDuUAb+p7SOKgHuKZyOJAwib9NS9/BHAFEwVAQjQVgnfVsS83BYrAJhZiESEaopWYg9+gSRnACMkA/c61SKlNNdISjc8G1ikrpCS/a9+v+7HxVKNK8LY/o/f/cQjP/3OW2++fufoDT19av/fffbxjc2uvrjIcfV/u9H1hp2WNQkvoSME6GTKSxZ+xZYWlqbKeIETjGuvce20Lq8iHnrRH9Lgg5cHV5Z9PjRUfPL5s08+f/Zff/LrRPyWm6763tdfe9vxq99447HXXrN10zXT7Tpe3gH8rTuP//qfPTJrMgICoQ5unQEzDAAKnRX78kLhUnVe3jJ1kw4MZAAq4vUhVY0MgdCFvf2i0H0Me6ed4dgG0vjSW/cdBct7vNuhL1roRhJdgoXvRohcmtx8Pbv4Wech3zlM4KFpaUMTjG6cm+I9g1hcN9KltlqyqFpW297ZObZzjJnNNKVMzEjs5iUeDVUzFWF2rTARkYEt5gsbfNeoWmBCQP9iKhLnwqz3bLepaRYRVTNjImZiZjVr2zbl7PvknIkoxFgGbV3UzoxDmG5tLZpGcjbRLqmil6qDgiY1QDi5t9h9vD123VPI9AO3vXZqiyjz7a0omlLT+Ek2BUmESIhMFJgDMxExEyGVydK0TVZlIh9bFSs1a5vGzJi5mkxNTLNKyhRCqKoaLAYGgqySpQ2BGY13JsxXvXjqpb3UvGv22T3a/qP/9kf+g//5cxvnwYgRI0aMGPEqwUhAjw1fs0QAACAASURBVBgxYsSIVymeeOLht731x//inheQIFRElrM0kbFiYoJSbNA6JgCyqYJm0YyaUDOBMCOCRWZ/EAxVFWI0NeIQqsgUkYgAOEYKEQAkZW0WZEaEaGhNm9pmMZ8hAhOD4WzevLh79i8//oVPfupLp87st2IKBM4ZGYAL5cBUdGtr67rj199x551vesObnjrx1PPPn9zZ3tne3iYkJKyqyg2Aq6qOMWqWlNrUpsl0EkNExCa1WQTAiJiZ3HSUiAIzArhnpXomsqn7ZhARc3BNVc4ZkZjJdWfbW1uigoDM7JbTiDipa6c5mEOMUURyTk3TppTyIs8ODprF4uLdZnGFN7sy6FXF0DEmw57W6aML4GXLZzs143AcvWS+S7qnpa1H5/qtZiiqhGCmqsVntpMtF+kd6GpFLnPj0/5P73H5o+xUfl9eaXCb9dc/9KV/9p/+2NE/8s8/8hU5gr3Ay8Na+4XCu3if5PUWV8SypeX+HVz1Pjm/DhuHlOKh4fbX0/rYwWFK/XKwzy9HQ31xsI0vAQBAVR977sxjz51djgphZxJfd9328Wu2br1+59Ybd97y2qtvO371JF6030uPKtD73v66j3zlO4NxlJuFuhVDVRFped1WAwydFQOWLX4vE/dvGQAR9I4aiLR6D57rPGNPsHZpDbCcG4M73eMOKLic0QYAoKLZsitndWBefG4MwlVG0JdRXa5W5Q+84NQ4woJiaiaSmnY2m21tTZkDM6ecVVP5igpB1Xn/5VGbGSLUk3roke0m3WDgZf16/p2WnujoHeYuetp9D1JKKaMQMxERYrHhXj0UM1PNfj04htSktmlEoJO6e+Pi50sBGrUk8pUnnkPTmtKbbty+YTvszRcgrUnxQimlfIEQCNylu2jmC+2NQD6xmqbxY69ihYSqCoSEZKImZlKIeDVDNANVyWaqpovkLiWEqlsVpQwLkq18EoL+2V0/8PN3/fWFL9KIESNGjBjxXcJIQI8YMWLEiFcj/uLjf3zqpRef+OjvK1hdVSBNFiHQyFwxMhqBofWsnz+aKaiAJtSMkKsQIgciqCJXMdYxcojEDAZADCFYymY5BAbIkpI2bW4W2rQhBmKE1mQxa2b7+/t7sa6r6Y5R/czJM1/++lOf/OyDDz70jVZAgVfsebGI7Ajpmquvffud73jzm79nWk8eeuihpmmuv/56JHQ1lo9azWKMTkC7s4aXCnQ5WFZtmqaqqqqKi/kCAGJV1SGaWbNoKLAhzOdzAGNiJHSWhIhcT+e1l0yVmIIrsstJKq6UIXDgIJKRKIaYJS8WTc4yn88X8/liPk8pnbeA20bSbYUKvkJsV0+srg7PSULsM6dfft9WXJuPQDDC2qF3qmoPOCCKCBb/jd5yw1QNpCsxt6zN5wGNIrq1AXfZ6w0R0Fb623ys5x/1JeBzjz5370PP/OSdrz/Kzl9+6sWPf/Xbl7X/I+IyXPnBmds4pYcs3qWf4576O8JulwWvHAd9bhw6XoP9RXr82TOPP3vGdcMAwEx33nztj33f8b/59tfdfN32JXTzI7ffeM/XXiw+Gx0L65UAwW9tXUavPNWh53/7F91dSdB5QA/rLfZmEYQrMYbhXmvLEA69N1Zr7q1y1tZx5usXy3XEORkgnSd7Y9nioD5kR9qW7ID13fEIHPSFYaCa2vbg4AAR6qoCpJxSzhJiiNQx9V1qgmqRMhNTYAbuyGJEomL5jMsyrdihv5RoYCzShfqQyDlqYhYA8O9T70llha83k5yREIl4UkMTGgBoGlMQLGVeTQehJwHIACeeO625PVYb3fGGyeR6SjlIZlBENAQ1BUM0QzBT8ViveUqLChgScYiRiMTjkGYLWjCzG3cAIbZgAmDAzDlnRGAmABFNCCIqTdMCARKZKlOoUPZFBXEySafa3bvugtELesSIESNGvGoxEtAjRowYMeJVh7/41F+gpNN7LyliZIDUZGnrKtQVM1pNWMdIbuPoZd1MVTIhYgyEgciILAasAlUVh0DEQKaoBpq1aZAQrUq7Z7VtmNlU2rbZ39sDwKqqbbojgPPFIi/2cztPWXaqiXK919iXHj7xwQ997PFvnpxn3FAZrqhh8eqrr7n99tt/9md+5sSJE4987ZEQQoiBiQ2MmXe2d1JOqgqIamamSDitplVVHRwcpJwCh+nWdDuEeYxghkiTunY2WUSYaDqZGIKoVCEQUogBi0pKidATfr1aoSIycxUrZ54NzIjBQvcoD4yV19Bz6nlvb+/06VNnz55NOV3oKi15mAGxtcbWwRVlu9YFgwBgaGsSaFzSwUdpbUgDFeKjI3nWt5etQ96qvAsdhxI4+On18lmIaCZg6KEIF0MjETN3yffFTdX56WWLbjs79Am4UBm43nXgKMd+jgY2iIt/40+/9N7bb9qqLvAPSDP4X//8wUvt+uXgMsy3VSJuSDov3+q2Ih4p1nH4HkEc3D998ARc+FqwscfLHFR4ZYHdQS3l3v7DYKgTBRH58rdOfflbp/75Rx/6kbce/y9+6vve+rqrL6qntx4/VuI8UlS1xGRqvrI5fWlO9cG6LUYZ69J/GdxyxTqTIlc9d7ZL5XVncNEdp3Ws9iAVAYGW0Smz7qhhaD2x8Tr36RS+PoAqECBd6DlODbpjBITeXgJws4HSMGnisE31URcTM5XcLuxsSjHGuq45hBgDIuScsiT2VdGouD93y50iMVOM0Y9XVMhF64Rg5VQbgKk6ka9QYgh+Nb18rm+p69r3d2spPyAntAfD5MjGRBwCl0UYDaxtGhNV0I5/9jEUcyQFOHl2fu/93+Q43d7auWl7wsgmLVURCQEUDAGIkUwF1QITOQfteS5qHpKMIYhqSqlpGkSq64otIKGpG3VASsmZetWMkIlEpG1Tu1i0QMSBEEC5WqSsGQw5ndl+6pq/Pp5uAXj6SJdpxIgRI0aMeMUxEtAjRowYMeLVhXvvvbfVhXCM1vLWNEDWPCfiSBgBGQFNtU2uTkIsLhyEiv5w31WcQmIjzGqSErYZNUuTpG1RhAkpsCzmKBkYJSfJqSLlWIVJ5LoiQxGJOLVpraHCuHV6v/nkZx+497MPfuXr3zqz1+S+5wEMgYirqrrzjjtvv/32l1566cyZM03TxCoyMSC0bVsyhZEMwdwx2CAwq+rB7EBVEVBUmkWTOJUn8ywGlnNumiaws9lBVLKIirpcmjpDyZwNEZk45ZRTBoQQAhgsmoWqBg4uB0spAQASgoGopJwPZrP9/f2zZ8/u7+23TQN2WeSzOPh5pdFxK8OeL773nsLoP2xrvMw56Ozl+SqlvwqzNSAxXL0oYEY9cdKp5oeuHR0ftjSsLb+XfPuFmSAbsJ6XhM1dnDw7+5cfe+SX3/+O83/4nq986+GnT19650fFFVHZX1SLl6S076bHancbWzq88WUf8JVKTTgybCOd3t0FBh5p6RjHzz36nfseP/kr77/z7/3Im4/ex+uvnQbQRZI+rFQUxf0tpWqgA1vkVazYIXdVDEXAAKlz1CEyVTNF4jUroM7B47Cdii0tV87R23A4PQvs1sm+2oOZCcCAy162P+wPEQkQg7sTl2SKy7OwXwCmBubfUGKqk+k0VlVvBVJK2ho4Ndxz66omkgfrqPWRPG/T9y91XLHEZgxMzahjkPuT4KfLXae9ssLagWP3w1SzGQDEECb1xMyaxcJUoXyxqvX1gQEE4CBJ286/8sRzk0A/dPvrbphSVMO2MVDt/lVCiATKYJOqCkwe4hVVMHQiXFUBwQCps9WSpnFbrc5gDERERBAErDVZEAMihsAGYKJqopKZ62nkpEhM757/6AEc/Nmv3Pbzv/mJK3h1R4wYMWLEiEvFSECPGDFixIhXFxQXlU0a2Q1V3NmaWpophYjorBwhmkgjiaxnNy0QTGIg9DxbRANT0EBZtG2SSgPSkOR2Pm/nTRU4EDECMwUmARMwYt45dhVPJhBrCFNTrEJFfBXGAFs7L5w6ePKxx3//T//yga+eOHMAhgxIsM4sAABMJpPrrrvune9854033vjAAw+0qY0xEhEhOYlcqjABGoCYuKo1cJjPZ2d3z1517KoQQk55Pp+bWV3XAKCiBta07WI+Dx1yziLCIRASFcIdEDGnrGqBOeWUcg7Mbuuxv7+vqnVdu/30wf4BIjKzmjZNczCfOQ4OZip56Xl7GfCKsM9DL9eXB+qS9HvYIGN82SHipvz4Vbiwz8zMnAFx/xMEQ+dKOmWziiCwu4d7V4RYlNCde+mGVP0LcZ922WygV8Tsv/fpR3/uB97w5pvOqUhts/zWR75yeXq+wKjW2DRbG+rlwEqbtnxxaad2OLy1FoYd4eH97fJooK94XsJ5YR35vvlAOnp08C4CIBjA//LhrybR//jH3nLEnhDgNTvxxMkWqISUVhwYzMTAQPGCrhMGoAaIRowqHqEyLWEp933qlssVhwfsm1495Yf7w67Y6ZKGpuFbyzNGXCTDitRJsc9/FpC5lEo1dba8H+RaHOJyhSWwVGcwA0RVbdqGQ2BmJPSCfP4l6MJwAxCRXq3cL29upiFZ3FfKWfecMxLFGEwLpa5maipOQBMxk5mJFLI+hNA1RQCHowEGZU3WLAIAhFhVUVXapjFEAENmUDBRVXN7GDHwwMWj3/xOnh1cv7MFNx07FkHbhWlyXyVAZARGqxhMc1VFJm6aVkSZAjEDWLNYcIxVXU8mEwAvFJxTSiklRmIKIXBOuW3bGNC0bRf7k+lkMt2qt7ZFNLVJpAVEDGQcgSoRmrdhp62z6Qd/6cc+8FufvhxXc8SIESNGjLicGAnoESNGjBjxKsI99/ypqiqfjcT1pBZpm8UcJFkITIgAKkqIIUQmYiJCItBAMInEBAggniZtSgakwIhAwcwkW11tTertwIGZmYgnNQdGVUMAIuLQMVoMpsCmRABB2nDf/Q9/6MP3fuPp07MWjJb2kAYGCITs7soA9KY3vel973tfTvnhRx5++ttPM5WaSyKSJTMzILgRc5F9ETqDLCIppZfkJUJSUwAAhIP53G03RASJArOotvP5bDZDxBDCZGtLRJqmUREOPJlOU9uaWQhBVHPOpur+kmAmIrP5rKprBDyYzYgwcBCVpmmcfW6aRp1MWS2TdUEMSJxNhEhHNBx6d8POh/XFh7YgdEaxyx42j+pwCvnhndYzzb3Uo2nng+Fbu+Tt3h+DmImwlxQCGOgyN7+k54OpCCI5+YKASAhZAQyJCtHsrtBeYsx6vwVTK+Ul14/gyCLol000DgmplWZU7R//8QO//Q9/8lzWJv/vZx5/7qXZ0bq4WJxfv3kltL3FuWDAOK/6FFycy4kN3CcOd3TBHi8XfUywNAN5JYBLvSl0ziL+zopDRXfTlrqe3V/FWuG3P/7Y33jb8VuvP6ol9M03HHv6TAvYFa/rBLOd54MBGKAhbFosYJBOoeUWpSpiHxlyvTaRAfsqYoDLGnpUeGqkznVazUOPK6Lv/oWnTfQ3tXZvFibaXEwtIoNP4lHW50GhwqIL7ine4aEe/mBJ0BlOEsON9PkyNAMA3QpWejQzhcV8piI7x45NJ9OqrhfzueRsABwCIGYvS+AmHEBlwURERKFsov3FqaoKOxft4bErgKi40lnNRNTtOHLO7m7Utq2KqIhPqmITjcVo38xEJIuICIGpalXXKkEkq4iZ9uuKOb+OAAatwMndxX0PPQb4lvfeedtOkClbZEw5iykxMEIgqKiUQpzN5jllQKzrmplTmxCRmENgEW3bNuckomDIxO4JguBuTmqWwFpEICLiiftoS05eupZjxfVWO188c3ovSZsawUAf/LX3feCffOyC02PEiBEjRox4JTES0CNGjBgx4tWCuz97t+WMrQhyrCOY5NwgIWHgwEyEiGAakAIzIbIXGwIkUDUBKaabBIhEjBgYGBmVjUiIkYhjJI4ESGBYRReiujNjIxmyghqimpoomfHZs7Mnvvn4Jz/9wOfuf/iF07NGQAsnYNblNTsXGGJ43ete/+Y3v/n48eMPPvjgUyeeOjg4iDHGEF26JSJVXRlAm1oAKESlIqFq5/br9QkBgHxgIqJdfUJCDsEVtUjEgTlGA1NTA6PAxAwAHIK5xzAYM2MIAOCFHFlVVBEJCau6clfKpm1n8/nBwUHTNpI7dmNpo3xhguPcBstrrBmubtzY1OF38dBHDnuTHpnJ3EQyHd7UEVTDdH0o9NCSlLbeULVQZqQmVvgJZzcMgToJZ9ei04uqxaq6EG0Aph0j1g0MB4wRwJKeOjLJegXpxQdOvPCRL33z/e9+w+G3Tu83v/uJR65c1xfioC8DDktDXxkc1j9vwmW8rC+Lr68CtVkvvN+FukVc5aDLLoMtVrySk+o9X332H/zEbUfsZ1pHDgxDiTGAGSpo4fixuwHL+zAkNvvgFDI5YV2WZVXckFpggKjgkUhwAlRMsKPR3XqjMOHlA8vMBhzYyh/WhftpKvEn7Ae2ee06tAXOfZX7Fs4x6dajK+eamOf4uBXVfk4ZDJoYYgjMrCL+hRjNkEhUDEBNcxL/6tbOjMXDcH6JnJkGMFPwOroAwEyIqKY5ZxWlUoDXvMTCYLmGnoD2HBfnoaETh4tozpJyDoSMEGMUIkRMpqbryQk+nmR2dpEf/fapnWPHrr/uurfefP21V20fm/CibbIkJ6AJjbs0lHo6qWoIwf/ZglVdAQACMrOqhsAilXYG0M41MzMT59SYVczT8g1hwacQUTQRUEEjzMrAERXVmEGqCLD/wbve9oG7ruhSPGLEiBEjRlwcRgJ6xIgRI0a8KvCZz3xooUlCBLJJVUlqZm1bBarqqmI3zUBCQDBCZARVBVWTDAhiuZnNwYQQQuAYq6qqAlMVQxUDSDKNSIgxQoxAAbJA24iIgfJ0KrNFczCbz+eihkjMBEjZyJAee+o7//rf/uH9X378qadPt2pqAKXSfe/y6cSBTafT97znvbfccsvzzz9/4sSJ55577qpjV/mzsWuuAQARPdU3xhi8NqI/Lee8RhzEKhKzuzwXlRNzCLFpmhjjVVddFWI0sNl8RkTT6XQymRBRzjnEiAApJdfKTSYTN4/emkyJaHt7G8qDNxThc9M0qZ0t5pfmZXs+rGSIH+aRX6XwjGx/vbRm1pWTY2YqimhLKR2hCRgIrIigIYZYlHW9dLGopjMzM5OqIgICqqqpGhh3VQsVzStslupsVgqhDb0YLoiXcdIv0MNv/vmD/973Hb9qWq1t/52PPTxrctf5+Ru56CmHYABrpglDM4fLM4dXbSDWBcsrNPFFF3k87PhQWtrU4xVVKA/Jx0vBL/7IbV9/5qX/7xsnj7Jz0Y92a8K643HPQZstZ7dP+l7vigiAX/zGC0cnoCtG8PJxZmAgXQlBW5qrW3c/duO09Zsd0R2e0cNIZSMdvrGK5YZz0+4aISYK6rkRJQLFiJ3Dz5Lwtu5VPyqCtXvXDXugMLFeinB9UXUl7xFPziXAuz9iWoyjV1tnyWfPnmnbdrpYAEBKaT6fT+qaQ8imSISIbcrdagcepaNO8EyI7GUGiQCgbVsP1lZVRUxNaiULALoI2szalBAgxti2bRaJMWIRrYMamCoiDh1TvEKvd+Q+J8W2xQSySW/e4vOYkJFU9SBbcybDo0/PZrvV33jvsa3pZBKzapbM5boamamJqoYQJ5PJdGt7f3+/aZu6qjrvLAwUmNnrJapATlkkm3uPIOScVZOae0eTKmTJOQuCgYhlyalpc24FADFCzkDSzOCa3TzbeplXfMSIESNGjLi8GAnoESNGjBjx3cf9998/a16awOxALFQTCgSApFwxhcBFJKyGoGQWGInQcgYRMAUiBGNCwhACVVVVV7GqIiECWOul5IFAVeZznR0wBxORtlUzDmGChgCxjsQoBgbEVU3VBMLks5/76098+otfeuibz7+wa2pec7BToSIh+ytCuva6a9/0pje9853vRMQHH3xwe3v7lptviTE6Wej8ORGqaMqpaisnoJnZDEw1p7TGesQqElHK2XSppzOASVUhUohBzUTFaWVm/zY3CrF8PMTADACBOTLXVWWiADCtJwqWc57NZ3u7u2d3d/f39uaLBdhFE2nnFYnigH0+NwV6SMQ3oKwLB1GEihu7Pz+3ipfuf7ykmTpx80rDxQRWTc0UELWonlcy840QAZz0UDArJgBEZuIVrYoIr7BRRkQ2EByqmYsBoZhIa9970dz3HN5q2bH+IAqTeem4AH380kHzf9z90K/97XcPNz71wt4ffuEbgzFcZmxqcYW9PQcueioMJI/rPGBvYLD24ogYEM1LXxrc3OMmme3m7S8Hl6iDnlbhv/+FH/rF37x73uYLdoGD4/Izhss7fa13K8pbg8Nn64WzR7F2KZg1qeSUOPXc+SkPutK13odpDz1UdHiBAACQ1vZxZbNqsTMmIr/9XcUL5TZFSaKoYEPlOC7jDX3CBa4PbKWbslDgIU+MjTPRXsaduKpEX/s93G3Q84bIhpmbkuQs8/mckIhpe3s7MHMI21Xl5H7KAlAIejfPZyRCWlLSooDIRJO67qxOCBFqnfiffR1C95XGUufAqASwC53tA3NrLI8X+gBUldBXZjIzVUk5LBYzmQuYllMOAGqK6ry4EJye50ef2fv0lx+dNbN33HbrhKTCXJE2qckpMZOBqVrgtk3tomklZxHJKVlX+VDNUmpNAYGY2JNecrOw2RwRVLKpKEhgJmJAVjVRMzM0QzVE5kA1W4s4YSKVvYUdvHhDiOmD/+VPfOB//+SlXv0RI0aMGDHiMmMkoEeMGDFixHcfi7S7VV/74n7DNYWKJbcMGhi95JKamQqYUZHHEQKgCYAwWGAMRBgnRBiYq8ghcGAyUxFJIkhF86sqmlvSrKoiyUopwBaRY8DAUQwzUJhuz5K9eOrMfV96+NP3feVbz55aLBIYkiuaukftYupLFGK4+eZb3v72dxw7duz06dN7u3vTyXRruiXFT7nk0hJxSokye0UmZiYiRDA1CWGNgA4xEBJRa2qIGGMEANVibQkAbU6myiGGEDgEyVlUjUxFzEveYUAEAnQDyrZpi9hWLae0t7t75syZ3d3dxXwuIufx0TgvzpF5DTBgn8/T8iYzjeWbeC556XlY6cuIXgQ3HCT2lQOLuWpHB3eVA5f7O1vhxBcRF+6oSBcNjIidTHJ+mZjAlZrOOPvFchZ7eSJ60nIT67lu6moXTY5eJP7gvid+/gff+Labr+u3/NMPf1n1Cvb4SuI8k/vy4hIJ4O9251Xk1123/as//87/8Q/vv4j+jnJOD+3TW2QcNBeh8J012ddVUwPTvlRp7yPcryPLleaQKbwTkwbg5hvdaNZnh7ObfazIFIGKsUahSoEA0Z2gYeg5cpgWBxsy1INVEAFcCI4AXcHGtau34dS9zMmFh14eWlVwfeNmdT2SqErTMFFdTybTGhFDjJPp1MBEhNn86xK67AIGr5JQTmPOmZA8nWiZgQSg6zR8V2UBrL+aTBS6lKPi+6xa4oKIxG6sBWbSjQHMLEpQ05SSSgkGl38EgBkCIgrCftJ0dvHA488IaDWtb752+4btACKaVVS1C1mLqrapbYVKSUxxuX+WrKJN2wIgE8cQmQMAimqWLCqR2QByFlEgAqDi/oTEZmCgAZgRicFSg6E6FmObdxeaQlO/NDl5111w112XeO1HjBgxYsSIy4uRgB4xYsSIEd9l3Hvvh3NuzqRnjDHGKpABKRt4ub7clqfFSMzEMYY6cMUooKAQ0CZ1VVdVFStCBDMUEUltagyKeYUbKsYqUKwQGMBA1QQhRCRCMFQxBRNUQwEAxSdOPP1nH/343ffc98gjJ1AtcBBRM+mz8w1ATAiYmXe2d9761re+693v+upXv3rqxVOTyURVc85N28SqCiGIiBkQlfzoqqq0Ky1IREwUOACvnBN/HkYsLIYT1uAGEabgzK4L59RANRCDWevOGwadqosMTURV1KmQ2Wymogez2QsvnjrY32+bhcolubgCDMjlV4amW+JKs3XOOxefUK8lCFYY6b50FRENypmBwdJa1EksRDAQlb4dKEYChAhM7MQEE6mKiAVmt3Nxd9RCwEBfBgy78MeG4ZbfayfHuncvPbpwoT0M/qc/+uv/6796n9do/OITz3/6a89eUl+XhqW08xxl/YZ7XmIHK9JkcOZwRZN72L/4gm2uXalDL8412ku90TrK8vJGI+rAAPB33vPmE8/v/j+feey8+y4Vz/2s7N9aZ3JLFAe71wiA4HcV0k1XX4SrwCx5KA4IAwDkLACF0ez6NCckl71v4J9BsiIiEfoCTsTW8Yo9iJEYVcuXjoeXnLNW9U8REefkccml00TpdrVPWI6vlBno/oCeQ8dV5nrpV786svN6QJ8fw/Z9zMscoA37Loe54ZCGBvpZJDCbWQghBO7HbKKAYOiGHOScPZj1pR1jiMQUQsidaRUzu7+Hdcyyn9oYQ2/sgr0DuHXBvG5B9+hs4ODu3mYmORmYW0t7KHeSJafcNHOBDCUC0cccDRQMsWF46oU50At1ReGOt+xMrhfNW/XWdgxtuwAzDsRMIrqYNeYFbIkIu/gAUagqLHOEzAANJltbopJz2ppOAaFpFm7RAQCIxBynW9umlpoWNBfzsUltzNlgEg/227wgfe6qR66a3QLw9CVNgBEjRowYMeIyYySgR4wYMWLEdxN33313lhRAFdKkqlib1AhYVjAwUzCiwIwIISAxMnVEH4XIGKqABIKWyYpUqhDOSODJ1CaAgOQeHQaWIbVmSgCQk6lI2+RWJCNQjfWO0dZDX338r+770j33fP7EiWfn8wUTITAgAfakQ6fPCnTDjTf88A//8PHXHT958uTe7t5isYDuSdi9R3MWM1UVVW3bFgBijF2acC7GDIjuxQHFE5JUJYu0besOG4tF48RmalspdAYTkoGpqKiU125taSZzZ0yICFXVmRdVwrjpnwAAIABJREFUTSkd7B/s7+/v7++lti1Ps9BrjY/CU6xzJXZoG1rPMC0pjCKS29wSDvbqt2LHnQ4rYZUTdhRSdZ0Y7HRtAB0TYkZEtCIxHoyop5KhEzx2xQURUbQYawAAAJULV8IGgx4BDcDQStdm0H+oPx7AkviPS2/ZQliDy/Q7/Wd/aH3XPQG77HOgli789RVk7L/2zEt/9MUnf+GHv0fV/rcPf/nKdXQhXLljXNMIb6T5LpqDvpgeh12sRxmO2t8558Cln7c6lrvpv/m57z+5O//YV85DcjlvuT6NL4T+XgBfFhHwnW+8/uiff+ZsQ4E9VcX9CpydtM7UoasLCMtfK90XUbOToYgIVOKCCC4+tX4f6IqPAhS7/xLHQkQ3oQY0wBAjRjB1+3h0dbVaVz0PzMlxNT1XPcGVsQ7WuH4R847F45SIHh47PzzlYmULHJ4zrv81JMJlcdZiMeQdw+oXSZH+LjvpfIQAUk4H+/uT6bQLIrm1tKqaJsGOvi8BArVe70xMHgZQNVVlFl+NRUTVYghmlnIKHIhwSIV34cLluVSVlBIRMedO8gyqggghFFcrDxdUda1g0CbJCUrF4H4dQAUAsbnZ86dnX370+a24ZQq33ni1qM1n84hGaDmJmiEhx8rF11YmNREhBiArFH021WymFlT8HC5yAoCsYAai1jRNzmJmcX+fiQEwN01qm6ZZABpyMKz25otZMmG65cUfPeDZP/ulO3/5tz5ygUkwYsSIESNGXHmMBPSIESNGjPiu4f777z+Y7S7mkOkg1iGQSjMHXJoPACIzBg4EyIgMRM6WKjBxYAgVSZNyyqSJ3SiZOnmSKZmgZQQDRZOUTUwSLOZghkyQs7RNmu+3jYowT67GHA5E7/vcA5/45BceeODrXpaoFQ2I/qQHANAxiGZ29dVXv/GNb3zXu9+1v7f/+GOPz2azlFPbtE4ugEHK4s+9IuLFABGxqmIIERFSStBRFf44DWCIFEJIqW3bNqUcQogxuuALEZtmISKIOJlMXUndtm3bNs42M5M/OTdN63wrIeYsKbUi/oiuL50+vb+/t8H84kg05Vq2+OaPWElx38A14WFeGGBATNEKLd2bYPTDcwnyEQjoDXw6gqvIoVjCqmk5Ra6bG5LQa2wUIq4INXu53cAtulizrulY2SXo5hrhXsVsoIWTKvI+E1Vnt71Vl1ljYfdxySZD4cysy+zuVJFLZe1G/vLK4bc+8pWfvOP1n3v0O489e+bK97b5uneHfHkOfa2VSyJ9j9r4xva7LUO19ZXDMoR0UcfoCmgAIMR/9IvvjUwf+dI3fcvqMeKhLUPged4zA6SlABoAf/7dNx9xeC8dtAetdEkM4Nyzh4D6W713X0YceMYPf7vjBZdN1L1wga513u5abuKBM3tfbRILQ21qplbFwIiq6uFBFRUUUGAiAFAzJkYCUSpq3n54G8/O2nkzMDA3EQbJAEBIPrbznysz0zUdOgyqI3rTXbnd4arceQzBCgcNPRG9KqAeEOiS00FK2mWQ+JhFxXlkYgIqX/SD2oxgZkzMzMTsySIuVVbRLKKqOJmY2WKxiCH04UaHmoqVxdMPQFWbtu1CG8U/BRAIKQRBBAMVEULkEIOCKooYoIB5sVkPKpCZiRkBnJ2lx791dhKfAcBJvbNNidNsO1JAA9CswoG3drZFsogYGhIQUfAYCYCqiWrOolk0KxgwMwXWWTlPhCQiBwezZrFoUwLAGGNd16lpZwcHZ86eAUTiGKpto6jIWG+RMdSvndgl5zmNGDFixIgRlxMjAT1ixIgRI75rmLf721tXCZykWE0C5Dyvohe7x1K4D8n8MQ2IEQmQAUy0zUKQM2puzKRFlQRqklWyaBG3mmYmqysOZAiSLad2kXIbiJwPADd3nM8CT+LkWKy3n3nxzJcf/fYn7v38Vx96QpXQ86jV1FQkOQ1inl4NqCbvec977rzz7U9+48mTJ0++eOrFnHNKKaVUKACArJJF+nxhTzfe29Oewg4hMnPx4mBaLBYAWNe1du6RItK2Ln9GKqJmQiQA8L4AIMbKqRDXXCPSdDr1B3dEqioEmO7v7+/vtwcHBymnoiy7DMANzJLhJlfTS4EVEsSIqKtMZaJ6RCHlYaY7WfJ2lxSUmXYK6BUCuuN8XfpotCIlNjMkBDPNJSObmBVgzf6410qriIk6LW9q2F0sInIduifuS3ED6Olm69SLrkfsKB4rCujCR2MZgjNW/mHEzicU4YJk/SEMGcONUtyVjQeL9Bt/+qUHT7xwkb1cGmzjtbeVd1/u5B62gp10d6ksLzdvv+XiOOLVoQ7bL9jQ48o+m8/AxcMGY7iUU1bFpW1QFegf/eJ7b73h2L+452FYnzn9NPVp3NOXvTJ15XD6ewwA3DS5u/X177znDbe99qojDu/Jk/uecQJaPIlWuyg/sOdLu8s4TMcAOFTnz98qiSulzGB/w67ss2xpSeamNqXOzZ+ItNMdJ8m+dApkA0QmVXVVMhJ2ph9rK+1mj3xBwc6uGnHD4rYBm948ZDNSrpOtjgOHemg/7v71OeMKvspR0yy8kGtdVYg4m82yCiLWkxoU27ZVMQQMgYkIAUVFctEFq6qqhhCIKeeMgES4aBqnlXPOa6y9LVlx7Mz6kZlVNYtY5+5tpgCYc4ZSClEJmYi0M74q9816hLWsx63BN549mzOQ8ffcdPWNO/zi88+x5a06hopFZfb0N13QDwhqIiahK5wI/cLitLta9w0iIpIlx1ARchb/otA2ZUSMIdR1DYDT6RSAgZgoxMkUQ8xISjw1yYH/1X/3/r//G39xnikwYsSIESNGvAIYCegRI0aMGPHdwd1/dXfW9NLB87HmremENaO1CEaoBEClvHtnHImdFg5ANVtOYIlRIQCDmUjbzFWyqVd8I2YOITIqmKa20bxIqQFCDoFCKESgGlHN1Xbcuhqrnf05ffWxxz98z2cffuzEqZd2tVdbOwtYag4VE+Brrrnmlltuuem1r005PXnixP7+nmphKA3AbUL8aRVVqUvcZjd/9ExjAyIMIVIH5pIFHEJADE5RuoUoc3AqwWsXeu06EXVv6BhjTzf0HTmpScROYS8Wi4ODg/lslnO+ghfVukf0o1BkQ6+K1d+lscKfkhNX0Kl/z6GuXm9qfZeBbM/dNKBTFyOgoeFKYbBO84iIhOpZ9ubTEaAEIQA0u6cGM7tibq1Hny3q4kEcVD/zq4uYwScsgJmamipzKZqphqbY0SZmnQJxObyhN4l1rEbhibDTex46rRdGcffAjjfs4yVdU8MGDQDOa7/wyuMKScA3apcvuaOjhFGW7Q96uuxq6Es8ijqu+NYjwn/2vre97eZr//GfPPDcS7PVZg9PmyMMC/tfCADf/4brfvX9dx7941988pTfq6bqiuUhrLcO2iQiXt3T13E/AOw/biJI5A4aSBt03AbWk9B9ZMiL45USeVZMk5wvNjNf8A0MjX09AAC0zqBpnYDedNgGLtv23xfae0N0qs+uKCvu4HMrS2TZG1Yuq3WBBlzduBmmqim189kBgFVVFavIFhCwp+ZdHVzWUQAiVDUVJ+OXWuw+JiSSzSDw0ld6ePy9LYkv/t6AlgCgISJ3a7WHObE7QgCXKkcE1NxqziZ5TSIOAAaoAGfn7bdO7lb8dDM7+J6bdqK0ExLCfM30WGRuFopIgSkwAbKhmqEBqPlMIEYGA1MDMP93gapklZxz5IqYTc0rGPtXeflXBJcAvQEDIMUq1FsCcNC0CwFhrRU++Cs//YHfvPsc12LEiBEjRox4JTAS0CNGjBgx4ruAj33sQyKphcgEcVJzQFKsIEoWcDPjbAAihlikz4pICKhoJtlyK7kxtkiBQzDFtklmRiGEqqrqup7U05rRcprtNQeL3Ka2bbauunrn2uuAmBEDYs4CGON0B3au28v87MNPfu7LT3zo7s+2CuJUoyoAqMmSeEMkohDC61/3+ve97317e3uPP/HE0898u6qqa6652tnenHOMkZkR0QvK+SE74UDEdV27JtofI6F7VDazENgMvIUQgldbEskxRs84rqo6hODlsFJKOecQQlXVekgfl3N2gdjBwcHsYHbmzNm93V3Juc9mv/ywixc+r9Efh0k5RE9ULww7ETEVKfHmrob54ctNZYBdCrb35Xn0S1p6WItsSEBjR0B36j8zCxyK0tgMEWMMCKAm60PpXDV6ExWgYgbAzITk5C4TiYqqCmLwWWGmilrcYwHBTJy3kk4MrsUgupBFRh0L0wk4cZAXf2QUUmegjS0RFQDQFXljIcRx2c+6BvI8tOblmYCHelxVDvvxbApGHKXZQsMbDtrE4UkdzqYBO3/kMfct9IPf2OP6/pcB2KmSu45w4wk8d9eGgBWvFk4FAIAffevxD/7qT//Lj3/t9z71qCgcOl2H3CSG2Rg4uP/LPPSoH/7kHa+76xfeVYVVFvm8+Pw3TmNvwoAdr9qz+G7QfGg4NuCml+sG9eehNKi9EXCxezrHpe/o7I5BRVgu1F0ZO69r2S8vvsKoQC+DVzMTsPMwuQOUOKgB0YU/spxchwZeqOS1HdBw0/4e+VJbmSiDsNXGHsAMCVVlPj8gwhB4Z3ubmFW1TW3KOcZYR88QUncqYiARzQBo5sUD3TQ/huAeU2bmPlTOKg/7k1K+t48Og5llER8gETFzYPbogKgiGhJ6uUAALHUoJpO2aVK7yI2p5D4iCABWTg0KwJl589CTz6fFgaZrv/fWG+IEUBc7O1vTqtqaREQKzNO6ipGJKYnkrLkr7RC5MlVVRYQQQwiVM/UiSlgqJboxV+lXrU0tIMaqRgoGJO5cQ0Ex7M/nL5zZi5JBW6Pqg7/ydz/wm79/vikxYsSIESNGXEmMBPSIESNGjHilce+994rOWVNCQA6padOsDZgIMkqLoISASITkdd0YkRAZwf+fVbIlQq2Yp5O6YubJZGu6BcQYGJmJiRFAG5Rc15MYSI/tqAlXVahqQIScrU1MEeMW1sdeeHH/oce/9cHf//PPfuGheV9RCTohGBh6GjQxIMYY3/Oe99x2+21VVb1w8oWTz5+88cYbJ5PaHZlzzilxVVW9RmmYC9zL3/xxt67r7tnSDTcwhOC2G96UP1GbaUrZTF3x5B8XyTm7u0PTNK0/l/Zkt+8mkpumPXvmzKlTp+bzmaogIRzm6F4uegrpiDTfUgW8vmXQwvCkAQLygPo5T1eIKzQWHGK8/N2+mODgQm9Exzh3RJLXIyPn5oyZbMm6rDfibBIzOyGSc5Ys7lQOgCKqoNQl8juDGTgAlnnSuxU4JwJeotAYiuHsyqnrhJal557ROipvtTrwwy/MDh9jz7ys/j632HKg5133nTgiEIYEmBtzrxCcq10Xgu3ijn+Vse5nT7lthhYSgyNAPB8Hfd3O5PT+Yu0YVhyDbXn9Vnq0QShgYP39coC9O/Hgmi2J5r7rTS86QhLtkAK6x7QKv/Szb/97P/qWP/rCk39w3zfOHDSlbVybPN2c9V5xeZRdhwiIr7l6+l//7B0/9fbXX9Qxfvv07LGTB94RFaLc1lXQxXJ+RSbc3TQGg0AODqyfywepeLVT6O7fTYGennMvNsMIoORfAUxEiKJONiox+UIUYgAANSViJgYANckih/I+uhGuzQgyUzUAP2pVPV/0ZfDOckFZmdaw3umGA6Ru4tKGW23gt3J47poVg5GU88FsBoSxqpm4nkyiatO2TMxEXUlAMDMRFVEiijFWsRIRUfHvPhGhkliCvWtTD3XXf1/DCwFdbufukMsA1VRFAY0ImRkMncv23VKMzSIsEFPT5NwOOGgzQOnE9guTk/uLp08f3Hb7m647fu11U6rJ2GSHOYZQhVAF8oW9rqOoNm3rgwkcsFv3iZmInXwHr/lpoKohxhiD1x9Ws8jBv1M8VyywF8tARbjq2DFiOL27v9catZOXwv5dd/3EXXd9cvN8GDFixIgRI64wRgJ6xIgRI0a80sjWBpomFSIKRLldgDQUjMmpXiQvoMfMHCIFJiYDJmAwAmDgSDFQrGOYTuuAxEhMDISA/lxuCKYipkaEIUyAt4AAVECziVlK1iYI3EjaP9j98tdOfOrzD37y0/d/67lTRmy6FMp1qdPl4f/YsWM33XTTnW+/84Ybbnj2mWfPnDmTUru1sx1C7BOrEcGJYKccmBncTtOMCEUs5+wH57aRPflYTDugK1hn6rnjAG7oaW7xLJJF0EnqnnHuCeheXpdSWiwWu2d3z549u7e760RP/6R95Gt1FJYQBz/P/aklr3Zoz3Nrlg//WQ5w7Qg2kEid/6kueb5Og0y+0QafPEyOrFi4DkeCgCvmF96hFqpzVfDZyxpdxO3sOR0mZczUPV4ICyPV5eZ7or7LJLvGluW8vJPlRe2PvR/6pdC8h3EuavWCst9zSizP+caFcOiDS53umlrzkpqH249f88vvf8e53l1hjQ+9NURg2qrCDVdNbj9+zVe/derXfu++DUM+z5a1d/uXL08HjRsVrJeE8+uRb7xq+g9/6o7/5Cfe+vnHvvO5R7/zma9/54Xd2bmHtX74deQfvu01P/POW37ibccDX4Tw2fGhB54B6C4JlfsSYe3i9YYR/YZOtj9cY1zaukHOi2AKVLxuCnXeB0HKax0sJMtPF4Jxpa1i4tG9cD8GBACQEnyAlWUQumyK1YmOqIhg5lkUUMJdm5XIK+diGQYDAKAu92KIDYsk4nJbmZrWr47WCaYH6916k27wIzmbKSJMRKrJNFDhi0UBDAihc2IpyyEiqJp4OT8RX0Cd6rcOqOZxAh+ns9KDs1doaP9W7JbVTjXdFb2ELuK1bIc8z2qi4iFh7Zr04ykBJgV4aZ6fPj0/8fzujTfe8MabbqY0w9yg5P+fvXeLteQ6z8T+y1q19z6nu9lNSjSpi0WJskeWZV0iR0Ykj0eGBzOThzzF47dxEgRwgAAJ8jDJWwA/5ClxkCABMhkDkwSDYIDIgGPEGVuyZNOWR5KtKyXRFnWhSKp5E/t+ztmXqrX+/8/Dv1ZV7X12d5+mmpQC1Efw9D61a69at1r71Pd/6/tnzA1TIMg55ywhNmKGFAABkdi581FDahjADcFAVZgZgJGQABGNiABRzAzIkIiDz0lTCSFcmB90bdt2eanHLx9uLqzu+W6aMGHChAkT7hcmAnrChAkTJryh+ORnP2lqrZ6EyBgCWiYTJppFagKiBQRFAI4UQoyxYSQ2QAM2JVAAibOmCYtmHokIVdEM1EAVumySVTokQCaSZCpmCs3Mn+4gtbA81pxMFQxza9dPTr730s0/+pPPfubffPmlV05UedbE1GURBfD0U4V6VjAzfeTRRz760Y++613vunHjxle/+tXYxHPnz282m9VqBZVWcF4YEZqmCSG6XUbXJTfWAHACmq3kkdOcxUxDCCE07psxek42p6r9I03TuCxaK51ZLTic/nYL0cJBr9frk+OTa1evbjYuvSx+1lAf5M8wVjuaux/hTETbw9tVtfJYCr1Lp+xaaiCeNiL1kvZVYEwu9c/zNfFXkTJv98RYCTjswS8Ult3RzMHAFFQAEJjBXEuPaZs5kixiBghMBAgpJdfQkYvsrSQfM98uDmhaYgxORvVZyxDrgJ4aSxw04Dvdeybs0Ovl2Ig0G1uVwEArbXlxwDaJVziwXuE6pqV+BAwuFv2glUv3XOAOcXd3vPPhC+98+KyZ7s6ITSe7h0amwQM9BwB9N+28Oxx47f22wz5vcZf9CO2qbP2D9YUNg3g7BfQYs8gf//m3fvzn32oGP7h6/PyV4+euHD935fjq0WbVplWXVq0Q4izyvAlvvrB4+IHFY28+/7Nvufizjz4wP0P5e7Fq8//9lcvaex952rqBQPSmujp4RwF9G8cITwW617tIAVDHSvZyISIAUBFEREMt1Km7FCEh5u0r9fe1xxTVbahy7qukuO0vX4nO03CxtY8l+1eJVYOP8cfH6wIiIdYNN9YnSDyz3r6u207YqnPQHhyra2aZ7ttLi4HH5pBQTfPxseRsAOuNipqoRo4MpCLep0ycRbqUYHtZYyxJXb2VWhL/Agf2FgVmCkzMHicW1TD4Xw3NNDOtIWFf/5moDh2Qh5PN0LCJ865NZq7u10JhlyYV/+iTBJevb/70r59q5vP3/cL754cPNNpauwxgESyAMWcOIoBoFom5aZgZR8L8lLqu60KIiChSepLAVCSJETM3kYmZWQ26nA0IgKw2BcGkW2cVRrCcsqS3X41tI//yn/6D3/ydPznbyE6YMGHChAn3ExMBPWHChAkT3jh86lOfgmQagTByjCaJWJmZgRgBTcEMy4MkqkpqN0mMAGcciAHJzLJkabO2azMVSdlUyaAJUXPS3DEZsRECqKiKqGEIhiQ5yWZpmxWYxdDMZgcZ4ZUrN//i33zxG3/z/R9eWYqYGaaUd7wjAQDAYoyPPPLoe97znve85z0vvvDiCy++0Mwas17OTG6d4Q+uTRMBUNVUFQDd/9c1ZVYsONhM23ZTnodFuy4RbXIWAPA0dK5odgLa9bDM3JfgCmjEYgadUgKAEIKo5JxT1x0fHx8dHXepO0Ui3NGb98eBMed7u7d6FF54i/IZKM/dttlWCb4Rfqu0nWtab8ALiNBv4lbfYb9d1Hh3ef2pYOx0jlXhMyA6t+w1V1H31nACOkNhopx6ECcviBC5xjMIeq20GTIPrho2qKx7uhKxCCmhF0rfC2HpKuxqtYC1P8YRgi0hZu2q8np3+/6Wh2y/0b1w0HeVT5+u3K5i1U5dsbywgRz/CZjtm3SKgAaA3eaX7tkx/Xj9sDWwfgS3u3SPFcmwh6IJ90AQI8I73nz+HW8+/ys/QoXPiP/zC8+vUvGyKKjU4GDTghA4wJ6lfg+Gu+t2Z9SgSvV6Lopal6YO+07I8wmCqiIRItjI22F8wS1yeHTZ8Wqmd50hdvtbBXrCtPwytncZYnVnwmgpLr9uxzkQR1G+3Xf7K/p6lbp2uYIQAocwjw0C+hj5ampmiDSfzU5/viegVZXqF0TTRI/QIREH5hBSSqrKbh1CyBxqEsLC77PT+lY2DPW7VWowmFylHpDPnzsfOSyXRyJpp6/8FwHciF05yU9+54VLT3z+gz/z2JsO4ubGqzOUhiEigKmqClgW7VLiGMm/FTxQ4et/3STlkWmvkf9p0X/dMTMAZDVREDNTUxVT8a0zCirUtOtWhI3l3Lw5ApmMOCZMmDBhwo8FEwE9YcKECRPeQDBARkbFOSNq1k0TuQlMZmRiYgiGCIRkACoiopaFgeLMDFHBVLqck+Uut5uckqQMasx0MF+YiWmOAVmMQE2zupdjZgNIbZc2G0ld4AihieHwxkl+5vKVL3z5qWeev3K8FmDWYqO8yweEEB544MLPv/e9j73jMUR87vnnXnrxJQ682WxEZDafI5GZdl2yklowAFjXdc4L55wQiZl63wxEVMVe4GYG1XdBEdEtLysB7U/BZQexVaMPB1ejz5QSIjZNk3Jq23Z5slwul5v1WuUU83X/+bg9suXXVpCZ3fWzZrsy5IF2PtW0MaUCCIS0Uz7BFiVtqiPGDUu6PwBygmRUPhLtkESIlVDFaj2sWhS4VIGoqKaKgMS9w0bho13G7s3jUAholEKmqmrZjd7btiCMnT6g+I64E6tL+P39exiOgdwvqmaoGdackBqLJne43f3UUj1eFL9219PvhtfwoR87B73u8t1OGVP8d2HrXh8M9Pc2VzlWY29hFn8S9/K/fHP9r77w/O4qUjS4qMUhuUqh9wQo9qici33HHTCE0Gp/lfWisNF9FRDA73LuU4ieLhi3B77+ssty3m1a26n7c4+X0ejXLSGw7gqub48dAvrUu+6ecefa1itnybJRm82YuYlRsyooIRpgVWdDbwk9qq2MHJ7Q3MKLyJP3+vLDHKiEcsvouMUzDkNU2tLz6DubYMhNPAzQwL9tCaHrNgYiqn3r+4oYmBicdPC9y1csfQ0EHn/kEq9vRdlElFlgBPOvnCTSdgn774icTZU5OBGfc/aNTUSeQcDttlSrA4n/kaAGWSWLmjoJXfJYIiHEA+CZgUBo2pVefVgeWJ5tbCdMmDBhwoT7iomAnjBhwoQJbxA++dlPggAyCiMBdpooADIgAiFYNlMlMMPCA5opqAaiSMyIoCKSu3Zt0kFOm9VSc2YgDkxMytDM5jEyaWYQApXcmhkT8ywiBxHbbFLq9ODwYrO4APHcM5/7yhf/9gd/89y1GyedEquhmKlTMNskxLlz59/xjnd+/OO/enx8/Ef/+o+Wy+Vms+5Su9m0qjqbz9UsZwFwkVTwpHPr9TqlJJIBIMbYNE3vUBljJCrKaERkjr3emYik+lqGEEREJDFzjDGEsFqtuq4DgNlsFmN07bNIbprGcx6ulquT5cnJ8XFO7kDyessot3CP1LPtshK4x3h0z8dyZdWxun7X8s6iob4vMDklnkQromkzc/duROLiM+qcjgIEJENKKZESMTkRZmbi9tDEIlnNQNQtSp0vMywiwbEX9LZ/Sc2ZaeZOC2P14701rZRXObdyzRHBU46OFI+2K3+uJ/upxb1jGKddJfVZa7ZDmvXJDHcVpCPC8F4tOF4PbCugccRx3QkjOX75YB3q+1m37Sr1l9kaoCHoU2cW3qMC+o1BFvuvf+9ry9XqdFQMEMFtkUUBAAhFGPTUErSPgN6OnNwGhIAoScG1tMSACGpgOqY0SyyGSHIGNWDaT84ibK3c+65+FnX/HVa/bQF0JeWrfNsJ6DMsp7ebi37X6eg0BKg36w4zPhJfIwAapE3LSDY/8HeZ2f1GPP2qh3XHVeq6rrd4tpqMt9pY+1KJSKn8HaEmIiEEAMw5iWi/dYmIssjY5ogQrS69RBSKBQeQGSEC2GIxQ9JNK6qAZuhM9XYHHS27712+eTh/un33o//Wux5tj5bL1dG5gzmCqmQKbIS7EzIZAAAgAElEQVRAlqUDsUDcrjep62LTNM0sNrHm3UVPjmhgkiVLVrWcUpc6AFCzLKqgBkBIhMSEnhuDkFUFGRrmTgFJ3/EqdAc8GXFMmDBhwoQ3HhMBPWHChAkT3gh8/vOfWEtKHJlwNp97rrXITRMwIrIZMaIymhIZ+yMUISFGCoGQENAyaBfJECKCHsxnloUAqYkcAzEZqGnOJqIS0FxUCohZNOV206YQFosLl3h24eXrJ08/891P/8UXv/DVb10/3nSiilRMfvEUcwHw7sff/ZGPfAQAbt68eXJywsyLg4OY43w+F9XKVheRsjtmOLncNA2Aa6KZfM+1gTs+u9ip6s7KFZumYWYzyDn7aYgEACklIoyxYSa39WDmXhDt8qi2bU9OTpYnJ6vl0p2FEemNFH/es/DZ7BRxuIeI2bN5vPzA08TQjoZ6iy6xEWlaodu2zuPzccS7qn/yzn1pVsTCZiZS0n9ZEf+ii6QRBM1NSs3IjKFKIotFR22yaqnawASZ86oDserS+aFWNlSkOiDfs91K2X5eS7PRa79qX+hW0bf3xrbRaI0P3idSeA/7PLzz4xY+99jjAQ1wqlf6gwWnxMj3blqyix3u+w4dNFzKdrcXlELunITwx4L/9c++880XbhExABjsVs9dFSAMmtY9BOv+guv8vn3vl60DRCOtMwKBGVm9hZHI3XzKskC3KRFPuU3jnrXrnifDaVONPpTksR2k/hCYAp7qwHv+NhmmmX+xWr/m36YkMwBVM0tdWq9WgSMTEzMT+UYUtV1n6iJpBygWHGaua/YVVcTAgJjcDqV326gO19YfcRtpVO2XYWfkTa23wy7yaTU1jczM1MyigmaVnDoVhe1BMQABaMV0k7/9wrWD+ezxtz1y6cJDi4sPRMhoWSUlSRzjwcHBar1WkRiinTtvqsT93yRkZjlLP119KxWgJxpQJDKwnLOUVIzU/8FBQAgEHDnMjWOnthFNIAwQlvET//gf/8bv/d49jumECRMmTJjw2jER0BMmTJgw4XXHJz7xiaMTvnBuLSnEGc1nkTAReCp3YLQAGIAJGEwJjBCYKcbQhBgDE6JKBkFQsEBEwIxwKCCKYBgbYEbQ9Wq5XncihmaKNouNW+52Oa267uhkdfHi4fmDi0rzZ1949g/+9Wf+8gvfeOa5l5OiIJsBUknQh3XDtJmFEA4ODn7uvT/3gQ984Omnn37lh6/MF/MYIjEBKBGJ6HK99gyB/tBLRJvNpuvSfD4PgZk5hKBqWbJvrVZVZmbmpolmKqIpCSKGwIvFgplzlj4bYdM0IYTj42MRYaYQDv250kVbMUZEVNXj4+PNerM8WS6XJ5v1BgqbiYZyryYM94jbK+DOgj3bz3dYFrTCQQ+cTM8PjPeqF+rZrHh0oIENWs7Cl+6wOObX21UC1qsgqvoFFHYcOPYqeJ21KQJC1/upCgB4FAEJkTxM4mLoSs6WIAS5etqvbeb2sKDaK50JzLRwJUiI2m+b391rv9Wie2ON/MJ3HL3BSNerOlJHl37ofQjqznof1zpYVTON+7Oo3QGD+tq1kmh9eryt06pM1+fOj92CY5NuZ8GxRQePfilHTnHQr6kpo76p9jBYLr7VnwAwnv8AgNuzpz8NDWz2E6aA/v0vv/Cv/voyxwhQbBJ2TjDVwVen3qSuzS8n9HGtvke8E3oKFQe57g55bWZQLIPLd0eZ9r4fYkxAq7qcdrgf6o3Ql7izccXAQGA8OmcEERkMS8zWcPZi5BoXHQcdYFd9X+t5lgk4uPPsLAhlhd6ODuFQ8qjncsonxyeLxcF8vghExMETJ4zXM3R5slqIgWCkgDYNboucM2JW1RgjEVtJ+op1c4lzzegO/UTsllaDHBudwhaoEmn/VnUvbw4cYzCEBlHN1mqqybYdolwArwBi9uL15flXbj1/Zfmmn33bo286p5tbJC1qd7JeNrPm0sVLJyfLnKVpmhhCYDbTttus2w1zENHNpvVEtTXual5hZuYQAUFERLOaAhIBUXVSMrEQIlJQoEzx1vL4xnKTNYerB+nC6u6jOWHChAkTJtw/TAT0hAkTJkx43TE74KObQvEQSaJxXl2fMRCIagLzLG0kpp5bh5kCM4IlohQCIRpoTh2ooAmTgYmppLZlxPlsRkREHGMEsEUzx4NDioFiIA5gCKIxdXORB94EMR6G5hzQfNPq88+/cutk0xkacu8qUIgLAyJijjl3jzzyU//wH/6jRx555IUXXrh8+fLR0VFsGhHJWRCBwdQ05wSYDYQ5VPWqEhlzcKuNrktZxMyaGBEJEDgwE7nZgvN9rp5WNdWcUkdEITAi5ZxT6tx/w1TRAA0YkUIAAATMKW8262tXr167du3mzZs5JwAAdRHsHbi3sxDEe80LsH+vHijsyYg0IdiRH46S/fV7rffU4E52CQPJ6Ym9ei6tkKyEzlCoKLGLzRWr6bMzF7tqUjCwsYXH9mZwRA6Fj9CcAICG9GKFtTEzzxjpBs2ARE5ncBBRVzG7+E5yMsGykdygiCUJVRQQkEjNQJytRgQkJlNVUW8FMdVGaJ8Zi5gAyNTV2eZC+K3OhMqZnB2VoSudhKfZ7aruHCnQt+mz/nK7Vx6pt2umr3vCmNipJdZL79K0lar+CbTguF1AqNe/A9R+tj7MYcMHX0Nz+llQiH8PB9SisdqtWGUDa01t+4LYdzgRBv4JUkD/4ZMv/fef+g7AEMI5fQ6H4LsPAAAJQwxlY8PolicED1sWlpkQPYyEhaaESlyeJqDruPY//H8slgzlpkU0Gt0xhdbsSe3iU1/qZYPfO9+uWX0F6ovaoP4WMFUraQ+xFFmiYm4WRAhkKlijr2X3xr7NQADjqENpRT8pekK99GcJ+tGY3j6l7rYqkQYYmWKbqUrerNemVrb7qHnWBGQij/QyqZqiBmIk5urLr2ZM5CMeREQFAYmZA89qAsPTSmpfeF3sjIQeAGQuqnBVFVVVYWImYiREQwQimi1scXBoeF2XS+kSVKk1lFCeAYAAIMALV27+4V88CUCL+bve1MQAmQAfvnQJEPJmc24+RyQRDYGZCZBic7A4mImqZFvM53XWYWD27yYfSiYuG2JMDYyI+1C3J4wozDWx8nw+Y9Wrx6u8fNu1uIqf+K2//xu/+5nbzqoJEyZMmDDhvmIioCdMmDBhwuuLT33uU2nVXThUQA3MKp3JGgzNxCS51EqJJCUVQURsmsLuqYmZIKjmlFpUJd9XbWqaQRUDEyEhEACasfPOgQ1RDLpNzlmky/P5bHZwSM18vcqvXrn14ivPPvmNb11+4ZXVuiVkBU8015OoViVy8ra3ve1973vf+3/h/Tdv3XzuueeOj49FtZnNrOuyZBEhZuIQYzQAQiZnRQ19DzgihhAQkVgDIiI0sQEAyLl4QKeMiMTAgcaSUVVzDlAk+xFmJwOw0qmD8nV5cnLt+rVrV68eHx93bTv0+5YG7TReGyc3oiTGXMh2Yc6g7l5sxGINp+0Wf3srh1HhNFIauvTZwJy0dbdM9v6qu6gBwKwIPweNoVN6ukVAlypg1etRoXDQTTjGCkUkAHCVeiWEgcg1ksTMgBkFmalkjgIDAKJQWRl1EkNJe8bFOUavNBMZkZJW5XswUyoiTEBAQsIySQQMkFCFhmlRKCg3r7kHohB9RsJIATvQNH2IYZDOVoJlLFHvOektkeNYNI2D9vIe5uGY9Sv+KNtzylnVKq0uUwCxKNB/jOiTEI4k+WOMm1GIyFNM805o4R6APjPLR8c0PQJa2UVQOeg+bOFBjYFJLZ831wM3IWTRnwQOWs3+t88+93987rnCqBq4O8G2E2/BDvNZhcFVK18iWYVNrqZJ1dLdPYXLvbVnZ8FdNhvsedN2X5mpqVdnzD4P98rtPf0HmfZ4kK0sKGXdRAJVH3J3cDIzIj/DhuAgApQv1d3+OxVSMttyPSpfT0OVRsE9gDrd/Le+zSb1szUxI5TREcsddpvNxlQ5BBFxPr8Mcy5nqhqRKLPHd81MxBlY86y9ACVLIFWS2rTsJtmB22gQUA1CsHeci47HYnlVMzCua+Z8caBZl13y8/rFrh9cAThep2fWV7/8N8/OGX/x8QcvcMeyXqggkapKFjBUtY4QwJJ0yECB3RBFFZsYiQgB63cOGpiKKEhdqlXVsqU+mYQ7dKFXkYNAZ8gHgZegZBRMlhH+p//s3/3P/+c/vt28mjBhwoQJE+4jJgJ6woQJEya8jnjiiSdSzvGgsWyhoa5dqaQ5m4iYZVRxuZeKdm2rIs1sRkgNB4SeOjMEMkIAYMBAREiMHJuDGKN7UJSHvKaBGEBzt9msT1aro5PVarNp259629sfXBxaXNw8ufrtb3//k5/57Be++PXLL/zQMDbMXTbd4sfQrZm7rn3/+9//0Y9+7MEHH3zxxRdfeuklVW1iE2MAMGstdR021MSGDrl/5HYPaHDBVElPj7NmjohEGEIQUbM2hoYIVQAR3KMj59y2rdVUSIjoaQxDCE3T5CxgwIiMDAhZsqq6ROv69euXL19er9c557Nukb6vOE2JYM0HtXPQX+iIgN75qNHd1aoIwL2Uz4vZvq7/JEJC6jdse7a/06Wp7ZIsnmnK+z/l7HueQyBXwAEAIbrqGQBEpFYC/biaIWDZys1KRTWJxOykjycrMzN3SVEzzznJXJSPIoIALoEzgC4lImxidEKkadDV9K4CBPfoIIwxOFclbm8qUrTSxHhqLO4EYmTuJbNWeLDSRifDsFDlAx1TCfsqqTUd03FjNgx6GegWtX0mICARFwpQB7ptdAnDSm1hFfO6qvSeLnTfsUmDf+tp4xYoC5gV6SxWqt2HoFrKmFWK8J4l0EjElfKvFGEf7gBAqKxc7VIiNHc32IoaQCVfISv8h//sL//Lf+8XPvCOB19Dh9wvHK3Tf/P/fOtz37sGTrIbGJgT0MyxP60G9hQAqNos+CoKBsTFit19jfwjRESBVVVytlRlrc5OMqnsJ6BfWyt8jpYxFlfg0hbZebZgDSLSvpCA32umBqjeOegGIP3HPLK7fQEP7N75ilYz/o0O+eyyvupQoxrOcuP2snDXPhOR5cmJLBaz2cxvCgMxsyzSphSYEalLuV+3sdcCVx04jr5qegK6t3U+fTkAYGZfZmMI4y8OROy/3/1+LO4dRPPZHERXJ0dWchjuhN9AATIYAnz5qe+eXL/20MEvPnIOOB0H1MWsOX94/uTkVkqZORpYl7vjk1sYcL6YNzESBVU6PDiYz+Yl3IkQQjArqnAfYRHJObXtxv9sUFXVLCIA/p1ICqjISQ1y4kybuR3bosG9DvUTJkyYMGHC/cdEQE+YMGHChNcRwhIlrHPH84jMIegizA8iNWTabdJ6xQRNCPP5HC8hAhBiDDEyq4iZEQKogAnN52gZNYNkAiU0Dqialier1WrVdR0YEBMzkmbNKXdd6hIYLkIM1qbVSbvsvvedZ77wpa9/6atPP/uDK8nIzJxvwP6JGNHMROzcufMPv/nNjzzy6MnJye///u8fHR23XSc5uzY1pSQipqoKIbQ5i0jOWVSVCMcEtD8Pu40vEYUQAEBEep7UyUeo5F3hRKqGN+fsj46ISL2iE9AzDnVdt1qujo6O1uu1SLai53pt0ub7Aqy6WBPJu2/Ux+YdRmsLhnucR3evAYjoO6Kh51wGTTgggqopQs34ZQCguJ+/sbGmGwB84FJGQjPLWQCACJnRKqOqAKAGIL2dAQCUQTdTURhU6mBqScXMQggGkHJ2AhoB8qATLBRTT+qaGWQRgKppw85ScZKlYv9tZpANwHyTeBYpn/X2MGGhuPcJQe8AM2eue0K0qooHmXH/H9ZeHaicKmzs5ZQjpSNUISHcjXS6Q+W06kJ7rTr2V8Fay8rk9lL2H+NNAQDQJhn4Z9wKmox+bodyqr957WOs3vT3pBovl0RXufY6aKc0Kw+NYxK/71W36bBh6CtJXf595tXj//RffOHX3vfoP/m77/6ZRy/cW53uB5741qv/3R89fWPZeR0zuMk+hBAAQU8TxC5k7kX06uwh9sbCHFjVNGfvbFUzNUSkpjEAU98cYyq658b6EQJ/fp9C1QD3N1d9G86+qhfn+K3SKylc62hqpgIugBZVJ4dH92V9uUcgfOdWgMdRsEY26kRHQLStMC+AGWr9IPmCgkA7euo+btBuNjnn+Ww2W8yb2azrOjWLMXhde5o4+xdqzk47k/9wVhpc7s2VgPY/MGgnnKOq3lkiAmBZ6oQx8+iypxd2cwsw8/0tvs+Fm+bim968PDnpNhsAAlAwqPlgAX3BJG5NXz1Zf/np77/rkfNvPhdkc+vCwfzRONtk2XQppU1sGg5scZFytzleHxwignRtWq27EILbdqmpiKiIiBATIiGYiGTJXdfFGJqmsRLdzN4Jnt/YxdoGUSWJhnNNpwD/4r/62H/8337unoZ7woQJEyZMeA2YCOgJEyZMmPB64dN/+WkD62ZdoMBNo6gBY9OEJlIDmk2165ihmTWLxSKGgICSxWVXaoYAhGSg6AkCzTwDPZiYaepMVLNKzjlLBgBStTaDdJY7yZmQQ2ioYcnp6NbRtVvdU099+wtf/Ma3v//CtRsnSKTmis7K64I//CKH+Mgjj/zSR37pwvkLV69effrppzmE8+cumIFITm2hjJkoJ3/g1ZxTzlkHVSYAgKq6VjcXMh1DjC4NduuGGGPOOXWdmhFRYGq71kxDiE5eq1MgBiEEBATtn9hxuVqeHJ/cOrrVdZ2q9tyCv/8GDzTUag07jndkbj2HMtp0bqeptLNICIsstOoZCRG5sL3Fl4Gq4K+K7wDq0Ayl1BcjTs6roGaqSGgAvkfb1Pn/oQpF/mbgPDUAEFIldsQAlJxOQkFTEVXzcRfJpoUUcR6h2He4Z2hVoTrvXK9lVdKnAGVrvlW1JgIQMYD5hCmd4GLDSnTaPXFjrl40NSK0rSSBRdholX+GgakaXlktoh4uAt/+9L6oe0fvSDDY3Q409JAqbuCiHfee6vC+Y90Vk4GBNB+mXZUel19h6KfKlJ6i1l/DDT5mumsZiDt3XP+2YeXN+sGr1caRq4ABfOaplz79zRc/8vjDv/HvPPZL737zG2PK8a2Xjv6Xz3znS8/dQECt9LGNto8YQn8H1SaZf6f0J1vNFzeS6lfe0vcWSAZAQEImEFWVcb/vOhn37hL3Cr9d1BNOmocirXwzDeGKM94yu60GHEd9sG+4gWGN5KgC7pR/1ht0HNoZRaHKnMGd3TElgjJaJ/wAEJgClpDW1rV9qVFNvqMIkWNsZkWJ7BJ1MGCO/Z4VKK75ZRdMCcIhmqpavyWlFO0bU8ZQRKubbMCMQ8DaOmKKIeacRAwJSQujjD7tAjMRB04p5+Tier9jrbDPYIBoREns+rr7+vdfSSrw0w+e47lws8kixBiiqUGI1DTzEFPapLTh0AAgZRMz6bKoegvatvNkxezSbwBRERVVQzUS9bH1kCgSgAKYMSibNbMGyMhQFdr5Cjb4z3/rw//J737lTKM+YcKECRMmvFZMBPSECRMmTHhd8Id/+Ie57cKsIaDm3CEHVGkDMCGAWM6dpUxgXB1ypUsqktoiKJacYwgHs5lKltR27Qo1MWgTCUwkpy6n0DTnLzzwpocvcAjACqnTbpNWJ9162W3aZnEA3HRGy1ZuXLv+vede/asvPfX5Lz617JIAMnCV5BZjAShkA104f/69733vr//6r3/2s5997rnnLl66SMgxNrGJXUrL1cpzIoUQVKU+7QbPGWgGvaKZmd0hZL1eiwiYzebz3pvC5VQi0sQIiGZqJszEgefzhY4A4AQ0mCesAwSEk+XJarVKKan2wucfM8/mRGp5WeTaA0PR7/EvLMTo4FYRdxPsIiATGZhrSgkpECl6qjAlQmJWUVOp2QgJwN1AdWCbB1Fh3ai9TSipGiLGGK04sI6MNVz+JmpgjCwiKlqdNkBScpUZYq9rBCTwGIn1EunAzhV4ikJEFNXKyCAYlLcQzcQMiKiMrsswzSRlJ6eyCphXGIqDh+85JzC//D2yvSV1lvqu/J5OHpSJRavtBsE4HAEcLHK3CuyHfKCl7TWwqM6njH81K27pw+ANIk4crveG+9LsYJPFitNBXzV/x7vCbegrvWxYZJMjJhIAhtvmXge0Z13d9KdM/xEl7QxZX/ogeh7ybkLlofsquFzX7/Evfv/qXz/z6oV5/LVfeOuvve/RDz32EN+j8v6MDfnys9f/r796/rNPXyk61mrjW4KHTsOJmJnsTMU6fXVkGeG7KHpIFkTkwJ4CNLcthUAcoU8JKNlDlLBvUr3GaWZmakVujEBMwGgpA6ARDZn9zniJHQU0ltkFakAlfOTrZrW0NnB1sMr2vNqSxd+h7qe3F+ztGWe8d48BQNn8c6fvLzP1EN1ms/FvkKaJTYy+nhNRjHNnrnPOOeeUEjONbKB8H5Kqmdt0QJ0kPb/cQ9Sjy+wnhKqtVhX/mt9sWhcdewzSrZOI+ODgwMxWq2VomjCbpba1Ort6f20DEDAFO+r026+sZoern3rkoZ9579+5NKPNzauLg0XgYGaARBxiCAailqj8lQI5JcmiarPZrGli23bJM2cQAqB5HlqwwMQhMDP4V5X6nyjIzGhAiE1skJvO6OhkfWO10c3henMtxNmdx3rChAkTJkz40TER0BMmTJgw4XUBRctrJd5QnOfNMQQkUJMkYBlgRkaaGCSo6iadrJcl0Y8oAgREJkNNqU1MGIIxNZLMJAkAYoDIiJGbOc8uYAzACCSmoGwQreHF7ALzuQdgdjDD0Gzsh8+8+Pmv/PnffPe543UrwK5chfJQ2MuHEQBms/kv//Lfff/73//q1StHJ8dqdu78eacSQ+DYxNl81kvtck5Zkqq60CpngUpTupKOiAwsRlYtzpKIZGYhRM8BpSpm0DQNgOacymZsIkQCM3HL0coUmKiBtW17dHTkxiOq25TB8PO+AM9S2kjmdsrmohccutayklxbXrRjWC9qBQAou+hrnKC/Xs65l/qqWfJfe0pPrff3HNw/y/UHPny4IgC6e6z2gjbuowhm1ueE1DH9WRlrzwqFhP60T8x+2RrVoDE/g9WktfppFLNsFSntrnyqd50WCarzvUMDykgjIReBHTM7z4hWHFuK6WoNBpwViNUzugxOYeC3N/FD9YsYHez/7UdqOOPUUPdc7L3ARiWPRND1353SrDBoeyjxNxrrVqBO7UH7CTDw8mWQ6zHveYVK6Pd34mtrSdkNUK5T+GbbKtKgn2nl2lsYloJeQVzqOTJMONqkP/jS83/wpecvnWt+5T2PfOixh97305feeungNdV5C9/74fET33r1T556+cXra0AKgcstZlsTa7g7EEo2OhjOwer/683AkRE5Vp8TMNOczRgBkNkAPIdbiZh4YInIl+Ji3Oz35qlw2u3I4iGQUxlYoH5KFIfkIRHoqMgzEdy07253ltms7IzwSaDFwmgQHe9+9PTl9pZ9+rR6T25Rzrtq6N3UoFYSXI5l031YxP9R1ZQSrFYAi9l8HjjknHOXcjaPCqsomJUEfdWOyUypbEkp8Tmo/W113wkOHQOmlrV4YfV+R+UbDKWIr4dYpqcstpSSxybdq3ppkDswyYRsoKpCCABueWIIoKI/ePX48DuvvvOtb7v0losXH3o4mETEJoQQIrJv6xGwbCoeATWbSZaUUgghxnhuMXOnr37yiGYzjSEAgMFgMILocx/ddCxwBIoLjLNmIXBVV2qHD2hO//t/8fH/6H/889NDPGHChAkTJtwv3H95woQJEyZMmPDEE5/oUjRmZJjNmk06WcxiQ4g5BZUGbBEDo5i2RKA5dW0bmJmYAAOzy45URCU1sxgjh8Bdt8ldMkOigBzUIDazxeF5RANUQNHcakomGjg280M7d1GbRYZw7dWbX/qrJ3/nf/hnf/ud524dtQbBdzmX51DT+hCOBwcHj77lLb/5H/yTB9/00NPf/vaLL754dHQ0n898l7driEJgfyZFhJRTzklEmIiIui4x02w2c1oDEVx15X7W9SrgCiYizjl5sfP5gRPQSKSqOecQIiHnnH0rcc5JRdEgpXTr6NbLL79848bN5XI5Mt+4V5xlp3zJArn/vS0fW3/KHZJWbW3NxnLE8Gx19YSBfQ60U3LpntbYYXyo7ptWVfdDZua6m15V9XSGLk+/hkSmqqJYkhViloyAIQY3+z7lFNrz6tTXxGXRxKMkV2p7rujmHtvsj7vKAlaObEfr6/RqdRKHogWWkldKFRGJ2Wl3K/wLgHuOQg21EJgamHHdgY4AgTAQzgItIh3OwsWD5vL1kxevrwZ5YmnpmN0dOOjCY+6VMxcmsOew97LA9qF3vgkBj9ftqs3rJClJVhUFEb9Reo7Uem5ul4mt+kk/7ZSmfieI0vsk1Dpv8WcDGddv068UsY1CJlsF1h+1ch4R6IsfndffG7WUGh2B3tYC6/tD+SVagzvN9pLcOdcJJiJCRmTCwNQEnkU+iHRuHjvRrz9/HUadNyLbxs0YwkI1bDO+yWsgpMwn6+tfz7Ke0x6KAnjTufmH3/Xg33nLxbc/dPi2Bw/ecumgCXdffG6t0/NXl8+8evLkc9e/dvnWzVUWU1NFAETuzWqg9yPveeTaHC3K72HqEu3exlYjeANvrao5ATEQUu9N7B1tgCWXKWoWs7JcmJlrXU9n+xzdNv1Nt5+k3o3P7KeRnSaGnUL6d/d+qv9gJdlhi2nGEvYzPUsmurOEJG3/V9JpUtr73r2OyjKisN0VOMzP/lsGkejw3OH84GC2mHddl7qkCs7JljKt5nhFdJMK/2rA4mplMMpGWMtEH1rP5TBen/1X37FUyhlY/rqAa+G4c84xRlU9OT7erJa5bZnQTEWzU9bFiweMDBqAhw8X//7f/9Avvfftj7/lEq5PoqZFjLP5IoTYpU4leWZBRCNmQjLTttsGLIIAACAASURBVO0AgAPPZnNEkCw1uyZJzmYaQnBzaGYm7FOaAiBIVhFDjIjBkDuFW6vlKzeOlt0mk0rKktaTEceECRMmTHj9MCmgJ0yYMGHCfcbnP/+JtoUmpiTahDlDmoMcUJgHYmZWYjM20ZxyThwQAEII/rDUZ9chImIK3DSRORCihRg5RObI3DBHYEZm4oBgQAooZuzp5xACQMydnpwcX7u1+cyf/uVn/uxz33n2peNVUqSab8kfc9VAmzgLHNou/ezPvefjf+/vHZ4/94PLP/jSl74UQmiamFLKOaeUY4whUErYdckfOHPOouJPuZIzc2iaiERd24poedwF659+57MZIuacuq5FQrcGRqO2XflDrJmlnNu2XcwPYmxS6gAAAFPqTI0Ab968eePGjRvXb2zazY/APr+hQNvPWuyhS9D5O3NSFYlwxEecUi8X6g2c7QWnmwygzz1oIoKK9Z3K825BAQmpCGixyt/cPbRkG2M2yzveqk6RlzyThDlnhGo8OrBge0bHJ4a7dpqZ7/oPMbjOPfcZKYnGnyYCbhgMUs6mlVuv9J9z1v0vVm1xkdBV4oAAiqAKZjpoQCELANjJpmdRwTluM0MrPxARTHdHEAEMq1y9Es2AY6oLiw7Rpe9WCdnhWmDwtWevOWfbK6r78bUiQK+U6Y5Ac1dP6YTujuXI6Wk3Ml+2PedYTx6PXVpGHKvHkKCX5feS5qrbHFhyRBh04qNtAlBo8ppbsL7sO6iw0+X0YuHrMkyfXX1/D9J0FDGQGiqo3h2IOFDYu0xxifKUq4z7yO8HhF4ljaVA6zusDJq7KtdWVIazOOr7q6vHm09+/cU/fvIFQPJb+uEL84fONYfz5mAWDmZh3jACdFk70Vur7srR+tWjzdFaODAzsy+zougMIGLXZlFFQqJCCPaMYc8PmqrnEvTYjN8i4vLYEsIxU+2pOVP12woRw3wuIp7tEhGBqnaYCpcHAEAIioP+entVGZI9Dpr9EsfwsRuvaTvU+Q7Gx2tUYO+Jw7VOF9h/sB+fIRrilLCb/OhdRdZnIaBxPwddIhh95GPwB7qn7zAzA5Fu0/rNrtZTzj4/faQIAHyZVVVV8VCuB7ZHIvhB/47Wr6PF86qeUKhn1xoXVrfE+Mqt7F/cPgP9NCI8PFxoarv1ygwIMXAQld4GygAVLBscbdo//6unuuXxwcfeN8+rJm+OJM3ni9l8DogpdV27AdDYxIPFgXes+oqTRHOGGoIBBEJSH0LNfkeYkJlmkT4ErgZqKJk8it9KtzHO3UazKaOkNfLhvYzGhAkTJkyYcG+4658REyZMmDBhwj3gt3/7t9/3vre/5S3nT04oMsaIJm0gbQI1jBGRXLenYiYGigTMFDjEEJgJFAgxVLURETAKgpopIAExh0jE6ImhCAAN2rVsluvNSU6diKgSYIM0h+bcS9eOvvbUdz/1mc//9Ze/8cOrNzddVkMosk3ofVZDiAeHhz/16KMf/sUPf+hDH3r++ee+//3vf+97zxwcLJqmGCP6w2oIHGPYtG3OGcy9IIxDUFFViTEy80jBiKICZswhBA4hhBAA0B9QoZo2qprv5zXzBHiqqkxcPTqcKlEVyV26fuP60a1bq9VKqpLrteKMCuh9FJ7/s6WA9iO9Ahp3+RQEOKWAHnO19ZCnWtRCnzJhnz8QBpYHrb9Mece7gqsCUc0MFMZ/5dwmQVgRphO5cYcLlr3/AUBFkJye3nEkqM23wgC6PBkJuTbKB4hw98LqZAGTz8OiXyaqHKM6ScW42zlU7hsvwF2hiy9HpSCKVNZUXdqJREgIooZgRK6AxkoBD7YlI42zE4lVkmiqYlI2gA8Cz+L1DAOBWdSoPctWRsZqgrhhKAYKtO/JvgB/v55fxatnnea7k25gj4cjI8/qrVrtFjWa3yNmfLsiPZtbnDJ6jfBWyT1d3HfLWCxdaGGqCuj+/y1av+8C12n2nYJV/YuVVO17wqpHDZRJglttKhQ3On88IiNLi3FohFXO0iql3DfB1azjosc3XJmSVtStNgQXvFjXI4/6SQdC0ItFImIOOWcV9d0MiJi67DcJYckyZ7Y1pFjX0iLSpqJb9oR1Axfc96fVO88MEInJpIZwSndZiQnVhtre5Rd7YxPcmiz9RYe4wV0yFu5M0IGkrQN36tI9EzmcduqU0aHxreK8rem4gNvgLAQ07Ceg+2vVqTsKomjlghXGmy+gvy0GBbS3k0MIMYZZE0IAxJSEmGMIpooGSKQlxkIi2cOEMHy+L2e05BWAqgICU/F48a8AJiqTs8yRQU1fJpv2k9eIiZkic7tZr1fL3HVgRghaLllvUjM2aADOMfzcOx765Q++4/GHDt88J2qXhETMbjOtJjVPAPnfCe4JA4g5JQAgZv87IotwTRtARL6byuoeLG8XAJqhKhLHEJtOkjaLk1ZaJaKg3KBtONhkxDFhwoQJE14nTAroCRMmTJhwP/HT73zLU09dfvDBD0TMjKDtirSLkS3ljEAxAjEguVsux5khUAjz+SI2MXBgREZy5RsiIqqljUlnIhgChWjk3ojZUA0ETGB5rb1x9da1V9erddvlJIjxMB5cDOceevbZlz/9qT/92pPfffnFKxRDIEziJAT40yghErEBLA4PPvyRX3z88ceT5K989asvXL68WCzatt20bepS0zQhhPV6HUKYz+dtu+m6LufsTsFNM/OHVxETkZS62WzGIZia+zNyCLNmZjPcbFoAICraVVXdbNZt28aSh9DMjImbJq7alYutCh/NnNpuebK8cfPGer2qBMPrHUU+TSLsZ3HrC60n0F3r5g/9tJOpDNEIse4ldytP52ZHbPNAQI9E0YSI1VzC6VNG1J7KoFOUuEOksnMugQNEBGJmYjOTnMEUjGi3ouXizJRFRYSC5wozZ4ABgBAMgHn3c4xk6KSgIWIIXGsiAECEKgpQvUDGVS024kROKwOoiIK5q7iYEiIhEpMamhayjBAVUQGVeSCgzXomqAp4rdj+uiCXANUUDE1Us3nNkAut7MzjaSLM5cA48DsDT+fmuXXse4uHknvNtYRVB10iOD4qI9XtgGr6gTCQSDamvnGg02Hr8zgW5NfZNNCoo7aU9wqfiFgpZuwZ4tJxWpWtpUmV5B11SyFU+zer7tL69yur27PSlcfEUWt6Yh/6sUMn2gid7ofKpVnNbmhmPU+MhYEadceImOvZ7+2mDKTkuDMrU92XMXoxPh9R1RAMENXUVMHDIsw2KtE/67QvByZEA1BxITIAADEhoZmJKvE4qmNmRsjIVFWw5gk5Qww6dJRZNdMvAS0cAmAIYIhWHaHLioAlfrKzCrroG4mqBXUdM6eAa/Sx3lrlLO+Bvne29Oinonx1gg67BUZBo22ieei+bYJ5q8Q6IccJA3YiatZr/29HHPflnDEctL8oF/NjX+eh8FM3oL9jduqyCGAq0pl1Oc0PDkIIKSUSNVXJZQdJH6BVFTCLTaMiKXWIVLMySh08x5YjR3HqN3NXpX67iZmlLnkouh9FN1/yDUlmQAQceD6bcQiL8+dWR0e567Iqh4CIJbtApeAzwEmGZ1650X35CD/w7tkjl+YiXXuSUkKk2MRmNosxptwulychRgBoNxtmRqLVcgmIMUYR6bpus9nMZk0InFKKMTZN03UdgBGxqhR23BdWwBBnoZllVOOV8gx5DhQioaExxn/5T//Bb/7On5xtoCdMmDBhwoR7wERAT5gwYcKE+4ZPfv6TJ9eOfvldbwWzEIO0S0YIgYlpPl/MQpiFGGMTYkAiDEQhAAAxx9iYZMsCqkTIaGhiKpI7SWvNCcxYGsySRNt2022WqtnyRvM6LW9pu2FEIzYyMDz3wKWHHn3HCz88ev65l5988rtXr90ysDZnrQ9hXltzzZ3mS5ceesc7H/vABz+wWq+/9vUns8gDFy8u5otyVmWa5vN5PTJrmlkIzBxcKuVKo16zycwiutlsEImJDg4OAgdT61IHAHHeSNkSC4wUOBiUXbo5ZzP1/cJm4E+hRJRSOlkub926lboOABC5KsVebw76TOhVrr3Cci9PscNIqORd39FtZkIkj+mvnrAgGHMWUH8DJXIayNVeRL2YGlxCNh79cgkFADCiYvTpAn0zQnLpqKkbWZxus9pQAXcOUauG4v6+gUnaHSIrSau0NgqHRHOIAkXIu0lpr/S3Fg9luoEVrlwzESGQ89o9XeKVAqfGzbnfUXf3t8JwLee7zExNQftt+aKi3XZ/w6BWHh/ti4RRjjgVABz234/4w1Hb/A2rnCEMDPPpnhju4v5y42sXAeSoUZVZtf516dCyKoy1uLVcG/fVDvqSKhespuNZOnRozR65Q6ZrdU0Ry+NaFQZ9qE2lyAdWrxL4VXTpE3RYEPowgEAprBe7j8odOOs97dsOL4zjCrBNpo7OGAWJhu6zIZpQSEYP7SCS1bAKIjIHb55lFQ+PuIpVzNWmKSeoZPG47QCgID6OWCTfZs53j2bXnnu/dvXQ4QhQGeqqxa7XAhy7JNcIooAVkTX4DbMzUbEyyVsTvg+O1NVjD0b3484NcPpeQLA7GDj3FyrlbO1auO1V9hV06sWdz99LQN8FNvInueNpBipgpjlhiBcvPBBjJKacUrH1xrJWum8GIpqq6JyJXckuImU7iTPOJRoxGnCf9IWbhp7AnTVN+UzpDLRqEm3m8mQgAiTyKoHZZrVqV2sdz8aawlMBEsDN1vIVeeblWw8/cP4D734c0iZtVqAaQpjNZqEJIrJerwHRTLsueSFy8RIgOL/cW39QtfYiIv86IqK+up6/t4kNMRth0qwcOCwQmnYjnUHWg8TZUvrnv/XhyQx6woQJEybcd0wE9IQJEyZMuG9AxXMPXSDg2XwOOQHkGc8axibAIvKMORIFImby1ENgHbvms+269Ua7jhBjIGOSnFQzgJhkFVU1pADISSxLkpxUk+VOcgfchPOz+WzBXaI2AYbzF98cDy4898J3v/XtZ1965fo6JUEUUdt6cK4sANHjj7/7gx/8IABcv379ypUrMcbmgQeaGF3ThEiiaqohBDMTEU9zj4gxNMxsBmrqBDRWRZWZLuYzyQIIi9mcmRGAmVQ0BFYOZgoIgXk2kyJVRXJiupfOOR8tIsfHx8vlcrPZ2J2YhnvCWYRse2jX0y9H1F+l1AANdhR2e3aNn1byGQCgVSsPs1NcYX+ZvoZjMsoIiz5ODRGMhpRTikNKsTGKgSi5+bgV9bJtMY+Ip7jzgaGAXjrn+slBx3daPFnL2+LCsNr1EiKgO4aDgYrsjNEWI2hDJxhrsXKpvi5Ys2T128a3KOORESxUPe94BPoOta3R7qWhQ2nb5PG4ENwlkcy8U3do4x3OelyO9affPship19UVrj/ZUSWurfEQG9bzwrbiFMtZG7fsjHJXrjc3rxit4vATk/10vSef64l9b+Xapr2KtZ+cox/jBjkQvRapb9Ri3l6X49ek9vrpnfut10CemCVRzT4Vjv2ENDjVu7UFnqPlt6noyi90UDBzAlorabn0NO+hVdWn61mCMyIIKJYiezx8NY6lauUm3F3ges55X7F6Lu5Vg18clslris32Y/UVnHOdIsPOCEbmOmuUc+efuoHYe+OjNM4Axt7F2yN5E6oafe8nWvfpkQanbD3nLs0rS5GW1GMrTt3TxVs9K/Vi6ukJJzC4qCJIYSQkNQ8oSsBIhF5Or6qQ/csrwBuHj0YBJXkrkNEs3wb+PFq0jKs8NsRRDMzY2b/88ANdRTMbcQW584BYs6imsczZNzOLtuR2PdfOn7kwdV7f/7ChfMPnMutpTYgxsgcSE0Xi7n3Us7Z51DJlNi73HgHDpPcI1b+lwX5aaICYE0zY2ZAa1NrgCHONMe0wOW6PekAFW+tr/3M5ZXddSAnTJgwYcKEe8REQE+YMGHChPuDJ574o2xmmfhgTvODQBrh3IygIYtsDWgwQUk5p65d57RRa9W6eWRU6zbtZrXSlA/n8xiIUJerY0CbzRvmxoy6JFlBFQHD7GBxcO7QwMxELZ2/+MD84BCIV8t1u24Xs7lZuHXcffHJp7/yzaezSjbIg9vACAjIFOPsI7/0kY997GOf/synX3n1hzHQ/MKhp9gq9omqDAQAgYtbQtPMVHW9XrsZLhIGJEIOHADAN+2GEGdNk1LqUqdZ5rPZ4uBAcm67brNeu6bPZYDEhExq5h6OZiCSVRUAmXm1Wt28eePkZLlcLrVI8HpC5Ed5PDwbr3F7EduIyqoP7WojeuD+12xEnOwnPmT7ZL39r7f7YH/Oa2oC/igj0jfpdhGGPVVCBACppIbJMDRyG97KwAB026d4fGZ/ZK+JCo5Iv701stGZ+66+O3cMtmjN8ZFRCbdryu1R9YV2mmEfjKrrb/XaA0dvY/q7HK72Mgiu0wW9TRt3gxyFN+77bZuzrtfs62ynu8IqCz50zk7j7zASe9+9zQk2EHCl405zUH7kDk4NBkDjAI714mI4RaeOSEXPqLYXIukODdlX3r2dczsa9a5v9VC4beV/AnCHRvTYu3bt/SBuL5N7S757ggHD0RTCUw77w81y54mMuUto665pAiETes7AEIKU8AExE3Hw3S2BGFxjDUqjwCEM1HOhmBGpBiLQuV0EUDURcXcOybnGO3C846TUssiNk6oeHBwScSfanRxLlr5t5TQDQmAANnj2pZPz52594Ci9+5FLD527YOsT1I5RAY2AYmicDXcPaET0FBT9pasPdd8E7I+4vltEEAMShhhiDIG5XZupxsiZJWtswkyOLHfd4cWHf/V3//jr//Z74EtP33UoJ0yYMGHChLNjCm1OmDBhwoT7gCee+ITCjCDaghcPXCIDApkFYhPSjNpFM9JsXWuSQDJaNuvMWjJFUDJ09+eIWB1rgQNRDIQBKApFU1BAmC3CbMZNA2SWO2jX8fCQmxkotpvUrtvNJv3N3373s5/78l/85Te+/cyLN47XSU1cCuriTQQEcpHy29/+07/6q7/2rscfZ6Yn/uKJzWZzeO7QRBGRiXMWEfHdtUgux1NVnc3mANB13egRFBBxFhsEzJIlCzEdHhx2XdelDgEChxgjAKiq5LzNHyMyiWmWXPx8JaeUVRURbty4ceXK1Vs3b7Sb9ix7k+8rzsiovsG1gjuSyT9G4I/IQb9R6GkjvOPY3a4hNvp5r589Xc7tzrynbrwDxXpfhmNvUffx1hgJVO9eyE/+BINT4ul9gunXUpB/9I1fcP5/jTOuls4a72xl2NvVO9N1L0l95pVwr2B9b6m3AVGYz+eLxWKxWHBsAFFUAQmJ/YvbAEQUrDjXu3/HbauDYAaeG3YkiDZEUNWchZk9Oy6cCrdWQ5zya5JkpgcHBwDQbjZHN262q5VpLu11ityAAQjKz7c+/MAvf/Bdv/KBn33fY49SezxnXTQEJmaiqk3TAMBms2HmGKNTzP4nClapvmuxa1vKPionoPstF0jIhESgOYEqEauYGnXQ3FpvXrm+PO5ybps3vXj5hYdtMuKYMGHChAn3EZMCesKECRMm/Kgws29+8wvXrr3QAS0wUu4kbZAAlBTUJIN0KoqSISc0JbBAQEgAASATcRObeTOLIYCqqQDqYh65CcAMhoAMcQ4GgAizORABmFpWMZWUlsftcqlJRGi9kcsvXfnCX3/9D/7fP3v5hydHyyTIgIZQ/UARwNlionMH5x577LGPfuyjL7/yyjefeurVV68gITPr/8feu/Vall3nYd8YY8619j5V1d0kJYayaJMiY7EpW2aMGKFs5MFGEARBHvSW1yBAnhIkQN7y2P8gQIIECBAgyEse7PhBMCxLdmLasS3bMq2LJV5EdpNUk93Nppp9qTrn7LXmHJc8jLn2OdU3Vlc3LxbXh0bV7l17r8u8rT2/8Y1vmIXn5g23JE2pNjU3a02JKO01RnoriIi0KxN5xLosIDLzLFQoIg09TqciJTO33T2AIuIRiGARC++quaVU1d577121f//VV197/TVd1wj/ieSeHkVe98M46U8yfgK76TbeJ0u+OTt8AJeBD6it3pZJ/wB74UfWoW+rQv0JH05vizcpnQOgRzWduIW3G6nxFh31jh+IR1FAv2mkPaL4+51U0o9+ae/3CRJh67rkU/pemQJY1wZmESmlMkb9QFXV3rY7jeFf8ZYxmUTtiDrTQ745bmZmUooIS9bG9dQd46Hsgc0aX00DTsSllFKKlEpSwh/yVsqQuG+t8CcPrn/ny9/46BN3f+bu8Y6sVgEngmfkOw2jrk+LiExmpVQ3a725BxHVWoZ9OfIWohRJ0jyPQkSZoBGZ4YWgcIqI6OThYCUFiZB7kNX+nY8G6sX76ZodO3bs2LHjTdgJ6B07duzY8X7xzW9+6Zd/+a/+/b//t0Q0+unqlVcERhJdeCqliNTCfV3hPk91krmIEAWRC8c0TXWeeTqkVeEwWSUnUwhhqugd7oisLxdoK9oSy7VeX67XD06X95e1rct6Oi0837vW8lu/97Xf/hdf/uPnXzMSFDH1dNLYNEdEzGAG86d/8c//4mef5iJf//rX/9UXv8jCTPy99RUm6k2vr0937945zAdiamvr2udpRu4qPTeezsQsIsJEIy2Xhac6tdYi4vLymphFODeKZlZKYaaAuzkAEcm6VdM0uXvrHYCZ9d5VdV3Xy8vL6+sr7d3jx6L5/bGQy/+2Y2+094THaKsfAiH7GIf8IFnQn4YBs8+Ln3z8wD569E580yffGkp4J+b6UT720Icjwk1bW4jo7r27AVZVCyfmefKaJsqA9nZ5+WArC5kENJVaHuKg0wiLeZ7nrpriYmw8tZuraimFhTevi/xxEQCkDKb7TECnJHo99VK4FDY3FnYX+EPm8XGrKMCy6AsvX37l688/WfQTP3v3TjWJpTCKMEsl4nB07QgQEQu7h6oiBs0dAQKzsGVNQqK0pY4IAkmRrLUL8tGqWacgIlIzXuaVp8vmK1USwcXPsPX//b//T/6r//E337Wvd+zYsWPHjkfFTkDv2LFjx473hS9+8X+7f/+lf/gPvxwRgMbSQi9LoUMpx0JTQREw43CcGCQitZTCQgwmYiEKuFNfWgDMXKeZCO6hrQHgotFbmDGRqZq20GbLtZ+uyRpTHI9HPS3L6eSndTn5S6/13/3Xf/T1Z19YujvDiUHMQggaBsrMQBwP84c+/OHPf/7zn/zkJ7/yla9+/9VXj8fjNE8AhbsQC/dbfDGYuZZap4mJilcAo+QcRtptvpwPh6w7hKzHtxWgP1sxupvHja+la3qb0tpa8s6ZMNtaa62ty3J5daldI0BvV0Bvx44fOt7dHOL94vHMJd5BFPzuhiLvgsdhnx/rRDt27Hg3PLprx+05SCB4eOvrgwcPpsPhcJiXdfVIvysKBzERUZ3qufAgsxBBRG4T0IFRtS/lz0ykqhhJTnCi/Aozb7VMb10UDY1/bC4caeGhXbMg4jzNhXkFTMmtI4PKhGF5TQBgwKr2wp98/+t36Kl7vzBPtfAUoWZhbu7qGfpOPXQEM4swESHcWjN199hacbsxgmf1DISbZx1CESJi7ZYHiYDDES0KH+YZCgUE7KWWCf/HM3/9v3zmH73XvtyxY8eOHTveip2A3rFjx44d7wvX14eLi2/0/qFaOXQ1Xwt8FjkUOlaZCjNRAHWuhQURwiRMwkwsIGrr0lpbWwsCSzkej0QUZm05hbswufZwF6G2Lm1dwtTWk7XlMNe79+7c+8hT2qwv2o1feeXqW996+ct/9PyLL78WxGruBJbKWTPMDUzMFIGnnnrq6aef/gt/4S9MdfrCP/zHy7J89KMfzX2amxNwUDscsuYPzLykAKlOzIQAi6QjZH7eTM0cwMWdC2Y2c5/n3B+ed6jhLMIPVVaLMFViZib3cwUhN7PW2vX19XI6teWUUqfM7/2Re0Dv+OkGPfz6hz763ofdxNnP4zEu8r2edp+Fj4d4K3W4Y8fjYpvsRMjaCar9weUbd+BPfehD7qqaThuOMAoSkYvjRYqaI2IQzETYbDfydT7KiaiUAiD9lMfjt4SZD8J3vJkx5oGtAuAY4MJMRF16hBNDmI3Zurk73EZFCuBWWVRywCm+9/rlN75Ln/qFj3/kQ/fu3LkT/RquEWxqBmOwwSnM3Jh5niYWydt3i4CHu4gUkSSXSylqSkSlVHczMwKkiIgsyxqOWotHWIS6TYdSDofr7qfVggoLLcf7S/+5Z5555plnnvlRdu+OHTt27PhTiZ2A3rFjx44dj49f+7Vfa+36dDrONQ7HuS+rUJlKnSt72NX1aeFRCSjMKYKZqshUqjBH2hOamZvBwExM/XSfmYWYPMJdzZiCCF2hHihTnY/TnbtMuPPkE/OdI47TRUxW7p5euf+V3/mX/+Cf/euX3njQgiIEYARc1SkIkcWIAjEfD7/4mc/86q/+6ssvv/ziiy92bdNcSylm2nuEBwLzYXryyXuttSw0nzcBAoGYiZjdfF21FOa5MObUQ5VSAzC1lBSZGfNWyWhTTJci8zRfn07rukapQUgbDwBmBuD6+qq1VXtf19UdQAQ58H5S/n+MlfF+OHn3j1/+7fGa4oftHvDYHfRDvrD44Q2bzZD97d5+Mx7pKuhNfz/Skd/mX3/0M+WnyZvip+ZGf4Lw6HkFH9TRPshefgcb8PFXZh/R8JIgmOlyur5PNB2O8zy31otwqSXciZi5AuFmqjYEywRmJuI0fS5F1rWpqqoSkYjM8zxsKxCZioS3OEdnYPisSnYgyxyHOwBLEw+Hq1pXd0f+t5U2HUshERCOWAOvriiv9T/81nefuHf8cx/7s9zrxDgcjta7dlVVYhIWMEW4u52pb1MzdwRqLbUWIiImZlY1IIQLsqXC88eMmkWA0xAtopmWUkqpPdii3L+8emPt84N7f3zvM0/pdz/ATt2xY8eOHT+12AnoHTt27Njx+BDxq6uL47FNhwNDk32LVAAAIABJREFUiYOZWdgDEQy4WbCbcMCCEBJEoIguzBRBboQoQoWFmMGABxcupTIo3N2cmYgRRJU4WAqIhbiU+eIotYDCuD5o+OZLr335Wy9/9Y//5HIxDw4CgSnc4UyEUU0opjo//fTTn/nMZz70oQ996Utf+va3v+1upQgRIkAEYoIHj+qCPFJ0CQBGESAnQng4KEBBBJGRB2tm7gHEOA5o0M9x1lCBsmohgYlQSqb7ZmMy87KcTqfl+vq6teZmo5V34fNj4O3FsI9HL/4o1L8/ZXi7Jn1bvvtt3vvhccQ/ljjNPrp2/FuC9xQK+gFfe6sY/rGtcCIitme09d6ur0HC83ycpymIMrLLAMKZCcwisRWcOHsgOwB3zof+mVOmzUwj5ynfelifTTAApBj5tgf0+WZoc/NwMwYxkQppJ7Xu5nHjmDHux4DF8f1r/dq3X/n4Rz/09J/7ubtSjlWm+UDT5GZrW5McFxECebhqi4hSiqmZG0ClcCkyDD4AMwuAKcsqwjf6292R2m9iB02mWV/RPJynSjB9cOX2C+vvX+rhf/pv/9P/7n/+e++9j3bs2LFjx44b7AT0jh07dux4TPzGb/xtdy/FmcHkrZ8CEcTqYe61SJ2OphbuAUy1lJu68mFAFZnmWZiEwRJEYCYCeJp4mrfyOAABTGBCrSDC0iCCUsIsekdvlw+uv/PdV/7l73/5y9946Xv31YmC4OEA584u3R5VDcDdizt/7a/+tU/9u59++eXvvfLK9+/ff3A4zFmlJ3NzkzI2s9PpemOQSc3M9Gwfmam7eStu7syFSERaa101IgLOxFmJfmyPAQABqGlX6717hAhLKUS0rkt+5LXXXvv+97//2muv37DPO3b82PBDdUyg93Hg985V7eYPO3b8sBFvFSy/S3rH7Tn5PtN0tgIJRGbqblyKlPLkE09dn5bTspRSmOBD75znIgIFwc1U1cyISFVrraUUYuqtq3YzGvlPOH8XW3UHJO07nu8EZhaWrHd8foITZ1Ce3Rxu4aY6ret0Ol31dTVT3NJTpxm0Bq6afuul15/79ivf/sSrH//QnamWSXWeahHupu5u7sRcp3qo9XRCRByPx/ONpPbZPcJ8FBjEMCrZflflJQcosjGYSKgIQYiEoX2ZnJ68czy9ccmnbrbUffHcsWPHjh3vGzsBvWPHjh07Hge//uu/DmrMFqROcrlcm661lFJLnafKhYgQcTgUIWJCYSkswsxMQsQUAhdymWepBHJqC0ypCNzRVxwOAMEU1rF2WPfew5RBxOxBl5fXy9J6sz/+zsu//4fP/tZvf+n5F19xgiGzYCNgQcQEoqSV6eMf//gv/cW/+Auf+tTV1dU//+f/Yl3XeZ4RlP+5ublHhCBrEHHv3T1KkVLKVOpwfHaLCAaXUoYLdLNmwSIRNLJckdQzzMPDs6gRDzE1ASQEGum6QQGPaGtbluX111+/vLx0sz8tds+3OYVHuaMPNsH7gxO0fpDX9YgKwcc71Hu4jh98NHrL+/HQXx/AKX5sB3kfB3v3u/+30U76Eb1QdjwK3n0A/Olr2IcSF+jWn+/0zs03bwuF3/Fj9E5NdqtAamzHQ2S2U2vr6brM08HNmAJhEeREgDNLKYWI3GNdl0xPqrUOFwszESmlhIe7d9VSkJroc+FhDHE0EVFrDQARmRoAZg6Cb5JqAvLRHyLhnnlhLFKn2rWYqnU9u0AjgraXHlgN33jhT/7JF//wb/wHv3y8ONjVctFVKE7Lkgz4svay9nmeUoitFmszVau1MjMcEXAnNwowgYIpIjzCA0BQBI34uDvgJBFkCMAZFI4AVZTicLMLJ4f+n//Nf/Rf/C//7zt0x44dO3bs2PGDsRPQO3bs2LHjcSBiZlOZ1zLdUVvgmObDYZqO8zTXWrimlHiukzAToogUZiZmpjTVgDe3FsJOFDCYRW8IQW9QzSJ/uiziStp8Ofl6gmqplYkjyE69nfTqWp/92jd//w/+6LlvvfTq5apAbq4234pUKgUB0zR94pOf/NznPre29vzzzz/33HNPPvnkPE2qrmrM3HvPbFT1yBpEquruqjoVL6UgDRfNzI1Abu4pivZIc+iUMwNQ7WZOBA8EIreLzJamkx4BICJUlYkZaMt6dXV5//6D+/cfrMua3pF/WvBeGb5H4W8e4ZiBh0mNxyB+3iTQe/SvvP/PPDo+wKP96A0oflzW5O8P7+KZ8RiD/Wag/pjwE9wJb9vMP1TX8/d7gB91Y/7A80UaQP3ATz3S0d5arvPNy+zbHudtyeXYRv+7fPFd2Ofz5+PhF8PoSntf6HR1WUspwhwRHu4RTFQKSqlEBHgaNDNz/k7INCkAgcgHNwG0XdWweHbPi057rt57Pt8zj4qIgrakpzSNJioRBMAjwtUteyN/EG3K79GONzpwQne89Oplif7n/uzPX1wcPnJRWrsmV1PlkZilIjJNU9p6Mcu6Nnc/zAcQJYHu4b5pooXZ3M09KCic4OSGMHgYxKkQSVpUiwiBQXLq0FVN1SXmiJVoN+LYsWPHjh3vBzsBvWPHjh073jN+4zf+NlFMU6/TfLx7XJvfOdy7mKe5CkfAPcynWufDLJTFeHzKfSAAd4RTeO+9tWs6OXl3W7w1144whAMkD+63db18cP+iCLsuV1fkLpyMtgiXw+GJAF2vp2e/8cIffPnZq94V0Hh4s0tgJjcLljsXF5/+9Kc/+9nP/p2/+3ef+8ZzzLScTuuymnm6PLt5KaWKLMsSEbXW3Ka2tl6ZI6iUkjWI1Lq7IcCy2T5GAJiPx5RKnU6n3jsAKYULj12rh0VWAHIpBUDvnZkJ0LXdf+ON1159zd3CA/D3nZL8k4Q3CWnfF8lDACEenaC/3Yzv6cQPf/GRyvH9hHTZj+AaflSs9w+gn358eFsO+vFahbZv/ujv9V0u+PEmzXs616Md+UfbKu/vbD8G9vkHnpIAf7Tb4kc653su7vpO//RBjbCH44vnFI1wXZbXe3/iyacu7tzNuoKtdyaapiilpkFWEseqCiCjy0CYqbkXKcw8TVOaOGe2U+/d3LNiYbLAZgYi4bTkQlaBAEFEzibRxEzuFFDV0+m6iAgzQMQMpjfdAYKIAYJ5PGj4zmv2B8++cJjkiac/cf+N1/V0eag1ws0sL0NE8nX+QcSH+ZiBc/OePzyEiYlZpKtq1kaGA0auFE4BRwEVkslN3ayUylJZynWj5qGImKY+YcH09LMvvTUMsWPHjh07djwidgJ6x44dO3a8N/z6r/96RHPv8zw/8cS9UqhgmolEO6yFG7tJgJWicQh5eNfWI4jAIgyKCG3dXSNMmBBqbUEkMR2BiPBl6UR07949RpgaRTkeL44Xd+Rw4AB1t9We/84L//hf/P7v/NELL7y6XLXoAaetqDxRAASKAHP5yEd+5vO/8isf+fDPfPOb37q+vq61TtNEIAKdK9qHRyqhaqnuTqA6VQIxZaVAdnNiFpbWGbhl/ohRyCctRgCET7UIRvGh7fgBNfXwfA3CPE1u3ltblmVd1/BApFiNH9mB4xF2gkQg3hThtKm7bjFf+eL2B7IFiQmUZiKbb+ZWTDEQYSnsPt9ditvPedAydui05S0/7HSJG3pxeINnQaQY7RlDh0VDiZbtwswyyjsysee9bF0weoHZN12biBCxu6upuW6kAYGImcbW3TyATLvOokxA2mVm7aYgBBOfz5EFoM6kYXZoKYVAHqNpAIgUypRn9/AopQTCzM5Su7MqMctjMgsxMXGMcEaM4Zk1siKKCIbtuAVQRQIRHjSuy/Nmb48cjyxyReFubsIyPNjfgtvZ5SCksj9vGhHmTkRF0nMmWBgxvsJMwqJmEdnmWV502LfnzZr5uRBn3mbmgXtEsi8REGGAuvbREebu5mHJ/pzZmZzXmXI/cseJhLmIeIRnMAkRAXWLCOIxDsM8j5Hm7NkRRBTjTpCXmtXMcoCMpWhMGPBWv+s8sN0GFZXGsGNEpAoyNhNYImHOlHxmzvWJiIkJQLj7dhaKEClEUPOcfHGrY85NmmtKDowkuUytlpKWrx5O2z2eC6m5e62VmNw83xQuqY/cpgmr5z/lwTHuZ1tOtxGZDTQGSq6WPr6I8CEaHWPPnUAsHB4ejhizOPxmwuYLM80Z5DEUqXmPaYiU05VH2940b5iXWtLf38wyjpgfBsM91LSUSswZ1YvwcV9byNDMhFlYsmXMdPMHHnPk3MURLszM4u4gKmnIcHZ+OM+h7RWBsj1ytEgpo5U2tS4TZ7+IyHlgExELm5qHM/FgGCWHF51HQQ5aMyMwiBHbYujmEdvQGB1ERPl+PnK2fxmL/JaKE4MMzWZRE+EcWnllW29FHjt7FkzYXCmY5dyqSbmO5cGDKA91IxwefUTZgDdtsrUiziNtu52HVyoP97hZj90jDOD80o0XRy4UZsuyEPPxeGQiAomwSHFX1Zx8kT7I7kZE01S3Zsnb8YhgMPOIIosIZ+9vFhwsQgAR3IMIGVoeKzMxiKSIkFDAzcJDWPIHhfBMByllbr1p76669XAgQAgCDLhW++ofv3Lv4uKTP/+xYzkc70mFCwUisrgibdWPt18zFEERUau4l1FbOZyQC9GUi23A3TrCwsxNPQQkzOJO7lykEAuYDrCDzBHRgjronsR//Pd+7w/+wz+Pf/p17NixY8eOHe8dOwG9Y8eOHTveG0h62MS8hBDg1pqYw7qFR2iBMZxBCDdyCMy1tSXcgkJYRAqBW2sEqqXwVJBOFcJMwkQRbta79XqYn3zqqd6tq9OduHPvqTt3n6J5DjW9vP7uN7/zB89+5zf+6e987fnvff9KO+AEEG5tmgEgAh/68Ic/9elP/+V/7y9fna6/8tU/Wtc2zwcRibTaYNk+OUiHqdbYSMNMbi2lZI1BIioipTIQ6RrpN3YZgx0AwDS7O5hyIzn2/QS1UZLRzUA0TdO6LO20rMvSWydCxMMb8Ufojbd7j970vyQSbgBIBB4414ra2FiAwh0EYhnukCLMQhCzDoC4YKMPtrs1Zqat9RAQkUGrAURUSxFhJt5qNwIYdEIky4PkJTMZmeCBzdQkuYHNqXOYaBMTb4QRs/BNSaXR+p4Vo0R8EKbCwgCZqZqamwiDGQAxiUipVXtXtUDUUkstbhsBzRIevXcgePCFkVRshihSC5+ELAhTnZJTGZ4sHrVWKRIBUzXzOlUAbkYED0/x+1bJagjl0nk8uaJAZFo1kqZ0r9OUNH1yJ+kJE+EERLib11pZJMXaZ29PdwfIzFpr0zQxc1ItyeSeidyNLUrqDObmbsw3VF3GY0zdtlMnrcwstZSu3dwA2hLeLUMcSdXp5mmeIQERMfXRdMgxHyKFgLWtdZoO86xqal21l1KSXMvJJSKOsDHp4nzYqdQzHQyEe3RTj2BhEWHQyC0IlCIRUFVmznBLUqLMg2uljYBOfmrwvwQmcg8zq6UIM4hMNT3iz/MsmzzJa9OeTLMUSXFlxi08MOzgN3b4zHiVTIxQTUuf8+V5Ore6ZT003iqh1VLcTLvWqTKzj5kWkhVQk4A2M7N5nplZVcMDoFJqaiQzYCOlqJnHxqkRY5BonqZJRGzbteY8jghiLiLpPHDmuzeqLgMYVERUzc3cTESEZQvqUE51DAI6aq0WrmYAePM0yI4uWxW49OAXEQRctU5TKYWJWtfeR3iJicBk7q33aZpYJJ2UIvw85EVKhLfWCkspUkpV7a01YWJhYenaA6hS1FS7IqKISCmmRkw1HxARILgPLvI8k241gptZKaXWmq2U61JOczP1nEpAcrgiIsKtNTNjzsu2XAOTdsc5EjDIRyYaTzEZHeFIFjKbgZmI8vbpHG4cQxXb8DvPrJIrhpqVDAJF8rPbgo+Nct+ec+fgDc4xWnd3pzEHPSKYWITdwzxuEdA4+05gKJEpw3V5SB9xOx/Pi/MSn8e1bPCIMDdz53CL8I29vYlWIaKtCxEOh7mUwoOhpYjI9s/JFIGAs5RSiltkLeIYj6KtEvHouOxcnMnfNOIYi+SITQ5/rYykyJjsHkTMPE3zmHTE03SIiNPpesFp1VP6h21RMQBwRPP4zvcuP3zv1edffvVTH3vqybsXYsskVOUcHRk/QnIAIai1nsdx13wOZsKWsJzjghHurql3VtPxSB7R4mBmEGcYzx0Mcbl4oy0ns//rf/jPPv78977wzF//G8/8o7f57bFjx44dO3a8K3YCeseOHTt2vAd84Qt/V82snNzjdLq+fP1V9nanllloLjRXSGEiwD3g6ZNspt7XWgXA2lbUqHU+Hg611KlOZRJKa47CJAQiaA/rwaBa5XiYNMIpwMwToaK7L/3yjat//tu/+//8sy/+7te/c712AzmlAuomnZ3AAZjFX/pLf+nf/yt/hUt58bvf/fpzz05TLVIcHghy6kM1OUCDJdx4F+apTswESuoqAn44zBHRexfhWiUizJLp4/NuMNVzpU4pf0uN3lQqAFUlKcn0tbVdX10tp6X3fuayz3ztY2AoRjEaYWw3mZ1ARFJKRBBQa83tpmwEh5sRca01W4GZRYpwyfTkUsrGGUTKt4pIgNwdCBpa16HPjAABpdZSCic952EWzEzCICJhYjbTM2fPzPNU4eFmppr9PTb2Poo7pTDWzKRIVrI8NxQXAaG3DoKwsHARllJaa9q7mmV5TBJS06Yqkp8SS3aG6awyzTEkLIjovWfsITbmzSy39KXUQqDW2lClUgpJBQQ366olIaLq2jUIRbhOdV1OXfvBfZrmaaoikiUrzczNfLiLEJikFGaOjQYVEUpiy8zM1IwRPLS6gxcuUkQqgHDvqswszG62ru36ejkeD0WKuyXrdnYwz6KdFKhTJaLeM1HbaFTHosheZnFzAHWa3CzpyxQsq5q7Z+I5E3kMdiapUhs8+OBrmNnUk9ZN6TRt+vr54mI+zMfDwd1678u6HueZidZ1jXBmnueDhbfeiUiESynZFvAhfq+1gMjd1SyALU0hiMjUQm0+HEQ4ImyT7iYZbzEUuyIU4b1rzkR35yJSSqbqm9lhPrCwmyEGVXrmnd1dexv8cgQN5vRmOnvAPHibpH4W+W4Ordm5Fh40AjMEcjM1U9MiRTZDgJTtJ10HBBPzOWIRY7gmWZYMaXJ3OXHAw1KgSgFgZiSc7N4m65TW1uvTqZZymA8Xdy5Op9Pae2o8mbltjvnMjEDvQ7rOTKqm2kupWXN2XVtvzXqfprnW2nq7vdC5eamFiFQ7C5OwbRw0aAuc1JrrUu+9936YZmEJz3gWJbGenvtnsjAiLDIaAVXL4gPJEprZnbt3mOh0unZ3YTlcHLXrui7MXIrUqVxdXYf7xcVFdrqcOciN383Aj5Syruu6tsxOwFhFKYdl0s054JMFTil6hgrcLSKmacpT1Fqzu9d1zbF3jn26e2ttnuf0d0q5q3D6QVHvCpDIiBkM32HmUsQ9TFVNM6q6uTR4RmWEpfd2Oi0s2XU1i9+WOqodJJdqdp653NamqvM8B6CmkmNOeDkt7j4fDtgCHvlcYBGMaGuGTiQX+Egv5kxwCe9dS5UM5IylLcNFRKZq7mOR8i3cGwiEu7lr3pSqmqlbR9LW2/DKpaC3djqdjoeLjPgGUOcpG3aQ5mN1pXMcJRfh7PItHhrMWUGQH3r03OQA3UxzIqq13uLbI49z+wNC4/bzCOvaYE4EkkLhmVDgyBgAXn79jX/1b75y9/i5j3zoScDrRBeHWqS4WeuNiZil1gJQBOVaRES9N2aaa6XNJDoHm6sRgYlUNSJGRAvDk4SZHZ7ZPPkXB6LeuXjjjZceXK5r+C/euVwFO3bs2LFjx3vHTkDv2LFjx45HxW/+5m9GeBFUIj5KX64bWS18mKa50FzpUHkuVJngIQQWAjxCJ1MpQiwzkiNhIiqlTrUkycXCmATCcIUQjFHE3fTBAzKngHB1xan7cuqn6/7KK2/8wZe+9rXnnr9/fdJgBweypvsNAnjiiSc+/vM//5mnP/PhD3/4j772tRdfelG1lyJGds7BJxBtyuX8lpoRoVAxN0cg4OkhkMpQ85EHPXjnoUfLjRyATYZ5VpbiTCudSVUAptZau3//jTfuv9Faiw+CfR5HeIsCOjXOYCYRRBABMsiqQX6J8DQNBW44gForsxD4/AHikQmexF8KwHMHi+SCxmdpyy5nKcKbQCygUkREAmBhFjEZrhpmab4RwsMkgrBJyQD2G5cPYq7MRGTu2pts0sgIAiiGmDgqFw+CafJ0qXX1CFfNOlRJc/ctS910qDKZOQB3YwSBaxEPV/V0xyDQ6G636E5bXzNRcjsQTxaJCa7aTJUZoAiYWhglA5YiPlVN94Ace6aWnFQq4NyyQWTQ9ID2ns4hyUFrV2aqRShFsmlMzlbEzmPPNDqGCevhMJ9T4909TOMGTqDC7OYZF0nnmU1MGODRvIM2NQelitZ8ywRn5hTGmntgaGmHv8RZAL9JBc2DwMyMzaciNX/MFO6tdyAJKHaPtIEYrWSbnwDBPVQ1iTrVPgpzqZ7z95N+yrkpwoggJjU138jfZIKYgygNQRBh3QJ+HkvYiojGRleNNoyQoVgfyf8ps0Va9gwBtaexTwzt/JClnrXb56z59IkFiMAIR3AQ0rmVkmgkEEE21XzORMq5zmTmAWeWFL0nVV2KdO0UKU3VTNKP0YxxHmkRoa5FKhGpG2KjWMMZuaZFb021uyqSOQ8Ot2TlUoPMhHDT7iJsailqzhCGp+k/wUwz1IHhxxBMXHNNCEdYeCRPjggfVB8KMyJUO4C0wohwtQgPFiGQdk3Z5jAp2UYaCCl7N1UqBZvJD/OwS2Ai8+jeZZVAMLGnaa47gYilj8WNPDDSEjY/ihzepuYBYg4iBDwig6k9a9kROyLMQs1sSKcBUnVVzTCedvPwXB/cAjQIX2xhrU2Qy0hXhkhrjwCndBgZ/wPgYQhkrBTh2keWQF7x2YFnXTUHQUaJpGTUlxicPhlukWMt8xa2O0bvDmKRapvL8ZmgTL8lt9i0zTlmsZk5MZgCOIcS85/cckLBLJjDeTQxmJGtHkHMTAiHRxCctrwd9yAEQQCiIJZcP8LJQZ4dDQoQ4OGqy+kkXKY6sUjqi/lmKmGMihFP3VKD+OxXMhTo25/ImFlsFjd4h6d2NsI2LuPmsIPbHV/M30KHw1EbTHWzJRnENQge8dpV+/Iff/9nPvLCVPiTP3tP1OK6Hw+HcO9tFZZSIiTTFAKgWqsIR4xw1Bg/I5/CA8ajAQjEpZRwg4cMhTSEhPOXWSCXfmO+d+/OZVs92nfvT5X0b/7Xf/0//1//0dv9ANmxY8eOHTveETsBvWPHjh07HhW1au/l4oIOF3eIfLHToRwPUu7UuQpqiUmoFjARAkWkDH45AAcJlVqOx2huTSNChLiwtRVhxBwkAMEC5uFOTv36en31+2QqiMJVu12f9LUHp++/vjz/0utf/fo3X/reKwhykN24TtzsA0uRj370o5//lV/5Mz//8bW1r371q5dXl9M8pSowBZsMSVFb2kZgo64y+TcyWTcCmaRPZBaq6h4iTAxP19XwTQy4XUScX6R40bYyQZq73BS1PXjw4PXXX3/w4AHe7Isab++t8Qh4O/Y6YuwjBzkQgLmTZJ67p9K71iojXX0wbpvQ8rZuK/+k20x6+sSmlvDMEiavGoAMrtBVtVIAoWYiUmpx99xlu3ZVNfeplCLFsn6jbanN20bdzEqRUoqZt7YuyzJNU5ECILXz2cqpK2Ti2Oxmhbm1ZmFmysKl1N5bqibneS6laG8gSrfW8FDVtBWudVqWU+/9cDgUESJqZ6G6j6TlUkraBWRjzNOcNGVrrWsPj1JqKbX3HuHEqVpF753XlYbKPln7Id8nYY9oraX4Om1AklolGi4Nw9KhiJUqTG7ee48t/T97IXWXqlpKnaZpnmYzzQiK33KETQaaiYuImwUiFd/uHhRn8+JBTEeKhVuqu8+tIZv7eXo3A8E8rCdiMw1InWZsviDMUqQMf4BBOYGYuyqWJTV5HqGt0a0RuK4t2V4arK5NdWKi1hqDmNl8OEKQ3IzGiJC8xBtHgjGUWeSh9ifqfY10hLARD5jUqmqO4d41qf+hmqQhUfdwN0+OPg3B00IBQK1VzVprtdasbHZ2n0h+mcatD1pcVdO2xzV5Th70p7u5GeAbpz++G0g1engGVrT3djgcYpqurq6IaJqmTLAYpBuRqqdZzbqNpckmAK21PHK6rLi5mC5ml5cPhqyVb4Zr9mSOf2bpvWcNtAxpbC4KkaptAKqniJhqTQvj9Dia57k3M7Pel+wQx1hRRSTbZ21rBjnSZODU12S/080gy72eF89zy+Twy5yJWmspI5mDha+2onOtNzdfT0spwsyt9ZzIh8PMwlfX10xMdNNfI6KYbt1M2aTC7F3TMqKUEoHeWgaixnTbtM90FNPeW++tTdNUSum9j7jOZj2RsvEI3NS4A7Gwe0vbi+0BpEnkA8TEpUiuACkVj8j4FpciPvS7fjgciHhZF2EuteSdEpFbAGYaqmamEchldm1tRG7G8uu1FBZer1eizEfR4fwuAmBZGm0RsuyRrOknRWLwwJqJLEzsZr11KQWB1nprLIVjcL8ID/MM2d5okLd0ARB4a9YY/H3mjJCkejdCARuOTxQevi5rlarTXETy8ZdmNrkU8DluaqkdHjZNaYO+BaLGGDsnc9web7djbLdG40bEA8Bmbi4csblPBbLGgDBfHI+n8PAwU7r1qCUggMvFrha7+9XnC9nPPPlLYXrq18u6Urj1xsS1lHk+dtP0b5mmaZomDw/zxSMzAJhFtZsphQ8rJHPK6KkqPERETc1MaiGWwLCLIUBtAfFTd47XrV+5S/PXL/6dZ5555plnnnmbXxw7duzYsWPHO2AnoHfs2LFjxyPhC1/4m4DeuWMihyfuHhl2Ue5F7xwhIDddtS/ewnNTytM8H48H4ihC6X8sJTJaAAAgAElEQVRApv3y0i3IaZ4mILStrh2upmj3F7VeAO1r76sU0XVZ7j+ohEJU0JgLERHk2W88/w/+vy8++/zLD5YgyFam6CHqlZk/9rGPfeYzT3/uc5979tnnnnvuud57eoZOdTpTe+FB4Ie4XiKUKatmMQkxpTszs9RSaw2zyV3jRqYUQuktOcqdFalmHuFUxcxNOzOJlFKgmtwctdavrq5ef/31ZVliM36+xT6f/3zvNHQEzG5/LyKzfyMpPRACsGTMUn1JlELus2wzeS+A3IbrsRdnSRZJR9MNp9eNc+n9eDiUWnrvyS6FB6uR9EFIuZsaM6+tMXMthTbBbN6uhzcWYcYt0wl3X9eVho9IirajrS11zb1djWZiZklltLn5WtYI773TyEavZqpmPDqK09/WzPq6llJEWNVUNY1Nw0NKSZV33k7vvWSCfGum5u7TNKW7RQpLS6nJyl0+uGTmOlXTpAK3qnqDQfHj8cjE67pm927Fo4Ycn0DpcZxZ+aWU1tYIMJOaAlFK0d7TejjvfSqV3iLBiy1tHIBIb61d8wmb6YGapUEBbcYNbm69SylFmHiUrAwOVeu9SboeZ+wiKICkyTZ33cjoRQ4PUyWCFClWVLM4IW1CvzSy6BFJ7dCQliJECjNntThsdd66Kqc7KVOWo4wIIibZyiMCbV0R4M1aVlXTCYTMPOLMTibNlFQ1AlKEidMyPkm0YeodbqZESIG/qa3rejgejofDuq5ra731w+EwRLuDV9U0uo2tj2utWXxPN5/ZJNTSvnzEdYbx9EBWw1vXVbV7eJ0mKYOdRyDXK2bu2k0z2WIMePgg55Lay6Y205ynyaGv65ps45lMVA8RESk5kZk5qep0LHG3dW0iMtW6LCdVa+sqtWQ2Q5rn1jrREJhfAyhlhItUN4fxcHM3tblO6QKMTdWZLHkpxdxOyylGxgPnwOQivjnqllKmaVLt6UpRawWhtZ668hHl2tyW00PAb8xeMkiGpM4zGENpI76xmVk30TzORkzuoWpddcvnGHG4/J+mg8evFczcuya1Z10paz+6RsDMwzWXIxAR2MNbU/dr9yCglAlg1UzJSBNnjqBMtclbWFXDPQnl9Jw5L+rusa4rDYbazzcFSof/cxRVlyVE0orKI4iJtKsCrXU1E5Zaq5mHW4dFjKXXzHtXtRtXqMS65tNquxDKh0kWYqWcFGaDJj6nAWk+UMaEzYcdZfpCKXWYYDQfVjIRgBPd1F+NLdxyE3TJwpKxmY+7W98ScW4so+nmJ0Eg3JdlCdDdO3eSOm/9xjeZeHh9mDtieEmdJdIZQhY55+ecL+ZsjzTAzGcP6BF0DpRS0ku/p5mVSI68rFYREflUAsAiUms+m3JR2iqbIgAHvvO9y6fuvP7Lv3j6+Q8f5zK/+N3vkuudw9xbI2Ce5xTdm6bLSkkFNYO2JU4Aj/BzXdczP05ngy0AGEL+CHBWIwTUPbgGEXojdz1OL9797M+2F7Bjx44dO3a8F+wE9I4dO3bseCRQUNAaOk8zQ9cILXCDw80cFBahbhpp/8qplRwbHQ9TtfDorQMsLBITwU1bZOmkzPLuvWFUB5pRmA/zHSnpfUskpfbr9YVvPPelZ7/9u1/+5vfut1UjIHTeayYHRwAgIp/61Kc+8YlPqOrLL3/3xRdfPB4PVYR4lJ3K8lkppNoYk0jCgUnIObmutH1IDbSa02BvkUUT02VSZBS+N/fcOOdn3G3bjTNtLrdm1rtdXV1dXl5eX1+/Sb73piZ/nH5KA+azwPX8JhAOt60EIYYMi1hSpmV+U+eKgFSAZ1FAZlIbJenORiKZRE9b2aVkeZhZTZNeLGYg8rFVT9lgY+KunYikFB4ElhJRgCJ8CGnDfSsCae7LuhBImEspKbVua2fm+TDnSYe0U9LsIiKilO7urfV0l6619K6qOs9TINwsbWfd3Lq2NFo1V9VM5I+ITZvM2Q1nZ+1knyMiBYbpmwFgng8R0buambAcj0d3080oI70RUmSv5gC0a/aMedpx8tnQNgV6XftWr0+TYPcwArIYprtPc5Y9jCVOyZbcImu2u8hj5vCjzQvFXTeJehL3hSUitPdaS/rMYmhIWU3b2kSGXwu20SPCqZdPirPW6axuTk4otZAAJT+6RQJKkvI5vCnpEeSELUTUTYd6OqsXZkI6tk8NZomIKe0+cjxTeobksLzxA6FzsUciMvdUrIf7xmKN0FXv3dyLFIzyhskwliSgW2u992VZeuu9d+29tyZF3CMAR5iZEJciDPJwU2ORIZ/cqChspsYZcclIAwDmkTeRWk3Vbp7W1WtSiuYegywWEem92ajJKanCTpsBbFRd1qxL2xYanGD65KRaX9zDPTaDaW6tISIdrkGoUpMAbb1xspOqbh7h3GWshG4RUUpLsXOaY4xaeYD2UdgwNhq0rZ0JkXLvjX9391oLMPS8BJIiEeFhoKFtz+PU0tIbnUBrV+ER/aIMYjFnZGsr7zmiYnRTDg4x6sDSNg4lbXDSa2GzQaHtKTBK8+VDJMe8Ry7sw/maRUo3IjKzHENuToDcFCv18/qbzkXnmnVJU86lpq56bWt6zaRI3NzGw4LgZuGR/iKpHc4jEmWQ0YSZhbUPW6FsX5ZhQJECbTMX4Uy76WpMtOVqRJKqdSsHmot2gMIj5cSj+KWfRxh8K5eaDbtVwxwV+cpW7SDXzCRwHdGGGX3OWXf3c+TJNwZfzc10KyE4XGBAcBsmNuN/PYiCIh20M0hMRHz28MGmVd8efNuDNEK1xymE6XA41Dr1vqgZai5Z6NotMtXm4QGRiTWmIoWzpq6nuw/SfwREm2cMmNnPi+Bw3N4c2CPS38ZlkNbncolMqVAWbL4rMVKgbgoqpmD69ev+7T+5/6VvvFDk4x//yN1uVEGliOkIGeay4m6gYKb0trrlTNbzrDIyuzZ3ILNMpHB3YuK8gLO/DzExjRKlXBEkcDX6pavfXstxr0a4Y8eOHTveE3YCeseOHTt2/GB84Qt/B94kgOJMdv3Gq0TK5N4N7hSoVYSpiJQylVKkztNUp6kyO0LdWl+v+7K0ZS0iU63rwhGm1il3w5TyIpyWRizTdHG4+8R8OE51hhSIgApY7r/w3d999p/83tdf+PYrpw4YOCnnTJPFWdRDKKV89rO/9Gf+zM996Utfevnl70XEPB+IORAyTEU1Ijy8q+VWOfdjhdLSgZk4BctSqpn1rs06gNxFF+FSazIadZrcvfe+tiEnJGYzW5br5LpjM5QFYKaXl5f379+/vLxMJhFvZp8fi3emN39rY70xzEMJ4WQ9LTUCxBhWmNg8X42YRMTNI4KTbY/YRFKNHj5FpBm0yNJaEqPXp5OqZbEpkVJU3D1lXwTItqvHxv9haPU2BwN4nWo9Cz+T0Yhofc2vSJcImIWpiYhvhE5XHenq7gQIszsDEeb5jqu13s2siHhYa+1IxyKFQClw3vRuBE4BaVhrSR9P01RrSWWfnYlUkd67byasRNwttOvptACotXQz39jxM4vBIvM0XV69oWaUenmQujGTMPXeQTTVyiIWqde74XGSTctvtd7N3TyykuTl5SUFpmlKG5OzArTITTlKIiaS7LZUu7u5qqX9embWE5O6DtoXJMzzXMM9+eIk5tJL1N2nmvJwzZTtaZqIOGWtRUStq3YzOxwOANZ1TRm4iKjaWZmeikIiEhZV9U20nhUiAaThukekISwCSfC5Owub2bq2WgoRazcRyQhTuGfhtdh8A2h4sAQIh3kGkGNGmITLclrW1uapBqCmRViKZLXGnM6nq+vLB8ZE7mGZp8+kN+rHtLaQqRRKDbh7+tgc5kmkXF9fE9E0TXne07LO85zKVtpU211Vu9ZauQgxXS9rREzTFBG6FW1j5hyBU61EFhGtdyGeSiGi3nVZllqLCKu59u5mFxcXZn66vs6yc6UWU/eATIVzGeyKDLcII+Cb6wgXQcD9KmnKi4vjsrRuGj6iRHZaNymoE1FO1STfzgrZ5BbbsoZ5lv0EkakRZXXGYeOT1gcRIaVwKW1tEZEOvGlunkUgmc8RDktitE6VRdw91MJDioDIN0JNavHNfSU2ZjLHnWUmSlYOpOTdmEcMkkWqj8Ckhg9d+7byR6Yr5LMmrSTCnVkoEO58dmDIOViHYc42DQcBvRZNxnk5LcnYPrx0E6W9PZEuTc1MrdTCZ48nAEAREZG2dlX1iPzAiMFE1Fr94Uqb53U7X+QwlpGhsomLMxtmdN/ooHzT1DJhIlTTm+LMiY+Y3DYhxl14FEFkaJMRg/QkD/L0/Kk1ww+TMAmSuc+UnGx2M3eLfLgIM4jCLN2DImw4RYkIUT5wXXPBuE1Ax4gxxFjCry6dgLt37/XeM7jS1tZ6V9W0pc8w9M1zcIurMQ9DHB8Fh5ExjFprbI2ZPxryp4WIICg82ta/RASijG3chruxj/qyt678nAk14uqBaMDL96/+6e9+9e7duz/3cz938cRHLlifujP1YwcwzZNHqFmb12mq0zSva9PWtPdS6tkQJr3s87g3bLmNcDwzQ8YCK1V67wFIKQBg3taF6gU5uYdi/fid6wdasWPHjh07djwyHtNicseOHTt2/PQgnnnmK7/0yZd/9iOk6+FYJsaxgGARlq6mQszERWiquR1EBJm7ezdb3Zp7pyxpFcMUmgilUC1sWeiJuEwzcTFzTAeeD4VYWJgrWMLhzb71/Iv/+vf+8G/937/2b770jRdevm+gAAdk6BChqeV194997GOfefozn//8X3WP3/qtf7YsSwSmqYI46yslh5X6TdXNnHFsp4d8T/uQcotIukAmZeObJ4Aw9a4RntTSKIkGpPIoKQyEE2XtqUj+bl3X+/ffuLq6XpZFVVPG9bbOzY8Gfsd/uWEfmUjOuq4UN529a5mZ0nXUA0DqEPP9FLjlRj/VbclV5ZZVMsWdKMWJZz3sdsazjyXcjIimWkZ5rK342za8cmeeRMFQid4yVLldkin3zFkVKtVwRMwyTFo9r4Q5q5dtbhqpNUMQ4Xg8qNrG0wkzn61sU2Gaos2U1XqEWwYnMMylEWm2ICJJ7CSnRURFSg6ANG8VEbN09dDj8Xg4HNJtFkOpCoBSQMdMtZZSyvX1lZkzc50nFjbb/MVTusucViFEbKoprc+SdKmUBMByQxgBSCow9ZJnXmjYWQSFe2uNmGuKwSPMtWxUpruBcJhm3uSN5t57n+pcpAxWnSnczV3VDoeZWXpvSUCba+9d1aapEpEl/8iU3gu3DBziLDNM9XoyhlsmfroX5BxkVXWztDrJPlNTVSulCHPYRp+Z5YBJtk67skhyi+pmEYfDARFLWq8wU5x9q8cRtpqH5yFKHp7l3TKgUksVYTB7clqmICostRTaDNC3cTEcJ4gGUZZr4jRNIiVdI3KibJEYgEDCQ5G6BWzSP97MksVP5s5UibkwFxbdyqHmBE9j92Fu4A73WipAXfuwq6nV3dWMt7Okq4lvFfBY2IdtCOfU0I2HHUYouFld+P9n712ebcuuMr/xmnPtfc5NpZJEAoGpRIChinJhHLgq7AamOm644WbRr7/BDXez56i/wk1HyA2HIxzhjsPgIizbMghDCT1AJQk9kCClVGbee87ea83xcOOba52TUgKOgGp5j4zIuPfcc/be6zXXWd/4xu87FECQYYpyz5ac0G3wNFRZBD0GU51H/BkOm4RrDxVkEQPUZVqqcWiYiDycabrCiQk2eanJj/bK9ID4mzugfAKpiycoPKKIVAQc92N6AMuJqa3XFTAQrEDpKcKi6sOLCoshKBd7t80qcmzjsKxOGEQl/nXuZBFg03FFE1HAHaz6FCawG2xxQ9IdioLGKlVVUVZRpYqqaUwKTs2cuX2I41hLM4LgB2eion30gbGXxBSiZFWKKvRWwDCQ8QgaFROrGe04ZpotLi1Ab+bJwCIse24CYl3Rr50TSsd/NLVj96gqBWKeCPmTu4o9beBUZL2BkD1xWXh53BfmXAbVFK1HRlAE0XET4WNCCpiU0/nutdc/LsxA7eNKm1mNzJhUEdXj/rifqIHeQ+wQeZy3O5QftnFikfCoIjOp4g/PNe2TR8/v90VECacx8iUBhhoD5xKyFvEzJUSL8uuL/ke/8rP/7B///K//4k9/8kU70WBKFe7NRrjvxxedSx++Xdfe+35nT2DHcJ64Y+JEfWzhwVOxx8lTNWN9cdtXEWGiNe3hul0iB9UQO/PwzN/+V//LX/t7yK1udatb3epWz+rmgL7VrW51q1v9LfWNt372H33xG+/+1mvUzZhze2ztBDGwm/RmJq2qVKUvtnuNPHP42NyvESPLe2tirWtLr4hkJuu2nMzdK4OJrHWxRqLUWomuL19FlloTtfC6vrx+6Ytf+t8/+7kvfOUbf/nuB4Ensyd/UE3lWFREPvWpT/2Hv/7rmfnd737v+9///ul0WpaTe7AkiSDLC+FUEXlgQ02tJpNRs8qHC56nCRrRoQUkXFrBtG1bRAx3KGi5IziOoLPKYEiulYBXXC7XV69erev296E+/41VVXNCelILmIWZak9YKuZp3lRVkeRiJlWFggFxk4XYQ0R6axA9IVXDSD5fcNcKRVqVTaWhcJTZRFP5SYCuipkadQyqQwAXUfHdMkxEREycUzDd8axwFqpYZm1jqmnNLCMinUiZD0FMVBTiclWJsKqYmdlkiUydGgJf5C4rTxVwjnXPgfcZ8YekODzZHwK0HFI98TyeVVUVIRpiJufzcnc+t6HhMzGLiYimjs9CvTVrRlQBSGjv1oyFw5FgmUwEXzlOyFDFiYsjastSVeGxz4hPxSTgFmSuXdyi6T0HFbRUWVX7sqAZszn13nEkPEZVzugqDJ5XikhvvVnb5bwiVa1SDfygmeyy/sRey56xN5s67rByt96oyEdMoyv0JiIChyHLwWlRJSERttbAzNmjBBnK7whv1oSlIie+tM2LdGrfHhDezdQjPKO3VlUsjDA0qgmkAYscXIu5nkxpmKASqSjS81hERa21okS6IBObKgTT8IiMyqkFV1WjBvUR12WnMmswjGclUyHHj4mGe1WxykHjxUR8ZIa7OyO5jkUgS/XWcAUSiTRtrc/mhFVrTUWu60pVpmrWMpOupCqmJmoeoe44ZWjXdp/sq8w4yr0ZmlVG88KAwq4641tVBAcRxs/ee+Y8k/FCvRtEUxy4ZsqTOMGF1QCtL5FiziIVwRstrYnw8KDMI6OSmT10riegrMzRBaGqqLLKajiUCviGioLSgbVERCKkigBHxqvCvMsiwqKi1NSFdtmbyAidp42pqkSV2ZAXp2bt6eTk2h24LEJM6TGvC2sT8i5zR2FHtw7YvMXRtAS1aR8TmXBtMkjPE+5cVROWINpEiyHI7pCMOrpQVMQlLAx7OCzGE5cvTMSiwkQlE+BRzAUkCqAoVBWTN3U69aiMcApG1xCpAFmz3QhWhorkhC7RZGzvn+RZzbbKpB1HYnnDmba7mKcLHrJtRGSENpsN5J1WnJk0b0ZoYYpw1rPL9tlboylJw8fj4+P9/X1r7cCCy26fn40fQYP2yQYO1pCIuGrCRDzverN5VlXEpCKuQVQ6Wyw/Oja0y+vP90Xx0VadHQacr0nPtgI3vxH13qP/6Tff6UL/4FM/+ebrr6l1yc04u6H1KbNxQqSmzayZ9d4NAjRWlbnmEfhXqurD04N247UIFUWks3AVxSizrtpE5PE6RNs90/uXy+OWzvlzX35nX75vdatb3epWt/pb6iZA3+pWt7rVrf6mqrff/nPK3/2tf7aI33/sTsclPNNXkWIq3y4UUTajh65XyoyMkbmJkKkQss64Wz9pW0i0VDi5mVoTbty6UwVlcCZVkhptl3j18t3vfDvdX9zdt2UZwT94f/2j/+cPPvt///5f/fBhDajPVZTFVQTBYuqq5/Pdz/zsz/zyL//yv/7ffu9rX/v66XTG01cEi044BtE03gJsABkaBtjIgF52MhOVKhpjEDGLEksRHNCl09dMeILd/W2HnZN2fdCYKgJOyYiIbVuvV2SCJeU+Zft3f3z7MQQHYeJ7Oh6V9NCgpyJNRFQFU+2xCQcCeAckULPgQ4A+cJw0p3TNbPfp5pGxhtCnbZ1wWOi8mbFL2vPdp6rLCvFXVT18IjsERmNhpv1pn2d4HXNvnYgj4zCTFWgJLPvHK1Ft1mAyFcG8O2i8LPIC4XhVZKYikrvic1BiYdBrBpErVmRFMmOXQkiARbS3bg19FJp9iEqwoSFmzI0T4pNYs23dMlPUVJSo1u0qzGbt1Bv2KgHxq+YD2WvVWuu9X9c1M0R10JbCy+kERWppHWZksEqWvgAdDFktIyOmD5QQQbWPhC9L660vp2XArpzZeleVMdx9ZDoRdDdtrbFIQuSd4IUnLyROJ+j7skNFVcVsCuUfOicFHNXCUD8ACDGzHBlCNlEhpLG15uHFNG3amT6GqvWlq6hHXK+X1joTXx+vVSmTvp2Xy+V8PrXWRHTb1og4n89ZNQJ0F9YZY8jMDFYrE3mEuzNPbrj7wLIAB6UII5ryer0S0fl8hhp7uVxll7Oz0ofHfBdSs90sn7V7QIkI1PhtDDivWzNTk71xRTuCwHc4zO4oJTVl5oxcujJRay2Gb+t6Pp2WZTmfz9fLZQyH27qolgWilDFTZC6LIZ2MWSB2ypSzd+n5aS5h/rWbVdY2Np4JnuQ+BWh0XZBMWHOwAS2JzEja/bo496sqwrOqWSuqjIQKX5UekREQ+4jZI2A5P52WCcL2AFaCVVkEvuzeG0IO3UONdZ/MwGHFNchCaEQBcrInbsImTyLCxJQTfauixyvcL/ewxwqzmjbDjEvEaaaJLsvJVIcPTM5QUZERLbOtSBOxzcy4uM53C9jTy2k2SKC7z94DU+TRGE3aOU7Y28iwPQLv5tU3Gy7wzs7oAQQ/Dh+Z2VuHwghwjaodcjrWyCMR1z1E5Hw6Dfdt25CsaGZm5hGXy6W11lvrvW9jGxsADjM4kVlaM3S5JhGbWXeMu0cg/bW1bmpYGbCTYxr+hefthkW4WcsMOi6ESDQORSiFaKYOzC5IPdFFnm54IlxkJBo5KveRmXq6RaIN9vj4uPQ+m0ZY8UWhygojEFSOiR/MSyGfE3fGeVbvRJS9ixlFpaIiE8GB3NPnq98hAc+xnvmj0/fNs18i4b6tW8WPdaeZkmgU/dV7ly9/491P/9m375f28bd+anzwjo9HGsStscoYV2ySX1dhNetTDc9ELOrcZpFl6VXlPlREjIcPUyxZXlxiKiB3VamaqFVRa/2FLtKUhd0vmct/8j/+0b/5T3+Z/o8//fHfQG51q1vd6la3+pG6CdC3utWtbnWrv6m+9Qs/9dbXvvvtT/+0dqMa2/pYYx00HWw8ODSyTauOOyK8qjc1PRCvLKokiJHrbVlYmnJxeeQ6xhZjjW2jCIb1y0dtV8pI9w/ef+98vv/hy8sff/kbX/rKN777l++v7rv3GQo0gejBKlR1Pp3+6X/8T/+9n/u57333u+/+8Ifbtp3PZ1hUkWVIO4lCVYUP6xZlIdIe86bQbOfIavQGifYYPcar9TYzl2qXI/eBVum9Q242FeEpUmfWq1cvHx4epvpch/pMfw8aNMa2J7hTiObrFZOIiSrrNMxNibho9/IKEWWmAikqU4AGM0GEc0/0ml8XPT4w7LHQkUWkWWPm4YOKhPj+7tDlhbgwhk/TsAm1d5n/rhN56hEejni4pyHrPQwwoufOhp7q+C6DRjhlHfbYw5S9LIaoNMiac/zfbNs2bOOU42VyLbATTG26FOHRJgJlhZimMuhOTGrSpeEdzaAQQee1NMxo0852EBhyCaPWxBCeiOh06pDe4FADQZioRE1V8L6iO8ChUkRMtTJFFdqKmgpziagKUe3OxDpC8HIO9c+/FpmpicgYAxFrqqLWiafdUlUy7TCPM5E1g4QRYxJvsau3bSUioIpxAmLP997MzEwx4a6mB2vbzFQUIuZuvoc5OqAgg46CDTezyEgqhUc1k08n9Hlaa5mJD0zES+8w0p5OJ3y9tckDgiSqqiTcackET2P6dqEnVpWKejgCBk0/rEAR4TuBRMDQ/fHJ8Wd8HghVNGEOYjt+ep5sRFnl7qZGzD7GdHruE/OQbKOAEuZEyhmRCH420UUYY+yqotLOu8DOhL/7qOOKwEVqzZgY4x3ocgCCjPULFwLvhBMVAW4lI7o37MCIOALSUCICQRl7G0ZytHPwsq01kUlQqSqzVjsXQlhEFXgRuL9FpPeldj81E3FrerdDVNxHDJGuqmbq7mF7fB5R5szVBDTJxwA4QFXHGIijRE03qwrC3eppVmQuazjcoxmA9thS5jbtydNoKsSn2mkwONw4z4kIpx8RubeIWE4nEnZ3nKXEFAliic0hi2dHjfa9l5mtKbOozs/M2GssRJJJiJScsq+JCDDlUQcLZVdpqwp9PjPDdTp84K7h7sJ8Pp/HGL0/mYJVNSLMBH/tzdBUFlHa2T5z8uO53RjgHBEV3cYWYVllagjZOy632lMRANhBA7u3RkQBOpZHZkxQ+zxJ9mM9T606Xs3mpZOVivuLhwDbX5k1e2C41oSKwsfj4yMRne/uEIvq7kkVVZNIpTNsUHfyOPZhxFxztjEwaHNMogwfaILGTh5n0YNU87y182x34SYd2BIRkp08Y61l5TEixVRyvADzlvTuw/UPv/jnXeVuaXd5vROHpTmJPEJNzSwjqJh5a62LSKIbWSVzfcKpzkSlrFTMJJmFlGXcuzOTkkyM51kqzNyUReW1u7uHdXu5jv/uv/ov/8FXvvO3/YJyq1vd6la3uhXRTYC+1a1udatb/Q312c9+5v0fXL/1n/9aZTWV9fLS14u4m7LxPvVKVBkqQgRmbjWV87KI8i6HqamNSJA6rZlYz7H62Hx7vF4ftut1XDeupEyKECpl6qd7Vn+8XGrQd99573N/+Fe+0EQAACAASURBVG+++o2/eP/l5jKZiEWURFlzfJyJ29LffPPN3/iN37Bmf/bVr756+VJE+tIxsCvMJELMWgXvnqkKC4aSq2iMrWjCbfmQaYkO2XS3hrUpnO1QV9i1InJsW07HN2fmtm2mcF1LZm3bdrlcL5fLM/LG35G+8VGuZ5nOLMz+Yv+rGe/BX1OizTJVNZN9E1prUxUtQjad8jO/Mu87RhS+MtkRHHiGbr03a0REl2IiU+u9QxAhokn33IHLtFtreadhCDOzWEVWx1tE5Bgb7SZB2sULeHunkkJcVR6RoZQ5LdPE02CYpWYq4hFzSyB6mmkmE/elR0yxZopPQHeIFnlk1I54kV3IS4qMikhRFtXeO0jPakYiCYe1qrUmLFW1jQ0bC9UyAh9S1BQHrzUD2qA1y8icGF+CLI8dDAHJmk3bvuihvHDRkXvWemciD5dda4aymTsIm3bT5LIsprau6xgjEkKwabPjnMe3IZYqM3agqFJROpsZJGYE0EHzjcyIoEyismbT2inCRMuyTKVs6mdCHLRLtPhOAMSryswQrkhEImqcRcVF7p7MvfcqCnwkE5ltIW7WoOEB/cF74UWIKMKFBRQdeCfVlIghHRKCzkJUpPWntLejmUHPJNGl9yIKd7BFmjU1bdaGjyoyYzRyIGMREcTiZkYsmTHGQPvEJuu5eFdscZIMd7wC7OGZaa0JzVZQVc0Lbb+IRNXd3T3Cl2WZA/WZRNR7h4P78nghprv7OyizV15NW++LZwCSkJH4w/RkRqpKU9u2EZM/bsTkY8DQHx5HZlpVBWfrTVWhts8dWERU4H2LDmBSVJWoJqaDqTUjssyUsYEmfD6fmWWM7bquSEU7LUtrPTOv18dco/eGBa1wPfAhIqPZKa21ypI5+6FgO8hU3FREImfWItZQnn2subCoqntkRjeFqr5uG0OOj2AmsxaZzGSt5eGaV+29i2IRIAUovKo1KyJtVlUifKD2h3tEmBoYxljKck87xBGJjP2KYeCS9y0QYa2syHIPKmbh1nTSS4gLgKPdQIuziJnNdFmWoorw5oZ/9+HE1MxUpbUWGbS3J7PSmqJ32JqpSGsmAte2YNKidiwVzl70unBjYKGMxFVI87eFmgANkJ5ERMWabdsId/QqaAepuzsTCZOq1M4sRrdgF+hrjJERO8inapLQiV2cnTnCfedizyQAoqrMy+WRmM53dzzJ7B450wl2fvokTVXREbAZHqfTSVXGPvkUe6IsjOfMHJFUE5q0O6Cfyc1Pf51/rJwgMPBfTFWIrTdPL5+tCQCm5/rNnFUP2/jS17/XTV5/sbz1RvvEvbhNnskIb2atNapCd6e3RVSrYsJRZpiuVCaLtNaUFZ1aIvw2Rawlmj6cipsSVRZJkhaDgLSR2l3TVw/K5d/6hz/1mX/yX/z2f/M///gvJLe61a1udatbPa+bAH2rW93qVrf6a4tTX755ItdmmrE+vnxPqay1fr47n07L8hQ6yJSUQelMiQfqHBnpRCnMKZoJnuSrurwS0ceHV9u4Ro0xtvAoaJIkLL2f7+7u7kj5rPY62/e+94Nvvf/tz3/5W3/x/Q+2JN+5iMxSNNGTVVUZb/38W//k137t42++8Zff+8uvf+PrmdR628bAg/HD5aIikIHwdFyRnuEeKsoilVEZxdW6+vDHh8f7u7ulL7vTNotCSBonVVXk8MGqmfX4+FhFIlyVDCc1ERWZGhN0N3YfDw+vEFL3jLwxd/P/x6PxEd/J/KGvMaQHhD8x5rNVoehN/MH0JNuUWjKTSbQZHOJZBdQwEyUlJylskpQiykxVAc0nIphThM2EiYUofWSV7JK0+6gqWIDB1BhjAGsAugUxV9IYA270YxMBEYXdjIjgqacimCupah3ONKD6MXNkMAubRKRXVhaUazWL68qH54wIwX1RVFnEleuG5gEcrH05bduUvWBJLWL38HAmtmatNZjuPbNZZ7FiWcd1Xdf7u3sWIa7ruqnZ3d0Z0JVMYmFiGREiar2Hu0ds7ryTmkEycY8xxsPjw935rrW2i2KJPZNVSLyEaVRIiAgMF1bLzG1sxKwqonZoJUUEirmKWrNIz4zKCk/hErHeQcMIIs4oAj1ABEIGkuGYOLPIi42EhZUZ2nQGyMnX6+MOUBa4EsfF0bKAzbmIPTKLKitiK5BGJu909nUOgzbciNMjmQX1TVUzKiIu44pDGRKQHqFFrtcVVwAEUCJC8hsRZSIOchyG68wcY4hO/DEaLLvDtKgoItZ1PdTYw0OKz7QsS1Y9PDwe+XLknDHWbY0IZlqWJSjXdQXnoVkjqutlhcAlLFUrhDsYZs+nMz4VMNOOdDhRU4Wsb7qpqaqt65qZrbXZyYm0Zr13CNA+fNsCkhk+6+PDVU21KRzQ2+YenpHC4prb5td1ZZW78xm4hnXdYC6GeTYzGP7u3tfhGZGVVlTFHjiie1Op0jMP0dx9xanbWtv8QugZEDEJe6iKiHiWuz88XkBKiaptxHAfDuwJZwYVpWddN163sYFYUu6Z5UQEmXg32MKyGgUCStXYBt6IiSMiMkRUJHBYcem13kxtumszjY2SsnIMr6rWGzFHpmcJlQiBT++ZkFDH8CoqEjFjlqgSNUQIZFWMOABH4TOuUyazQzLKRwhB3J/xjNf1iuuo996sNW6ENoPo4A0EJJqiZaiodTVRrK9VkelV1FoTlsfHS2aJChqPrS0A7Yg4iOK0u+aZMyPWWFVUJzrDw0OaSqnsLVWTRkJRNbbBxNbNTMdwnJPMbIZeZSVi+HZruTC7x9EWEhUhht0Yl6ivG2cp848Qe1SVqnAPnQ0EPgz+WHBIVagyY891FCHC3IYwCbqK9XSPPBqiVBnr9frDd9+9u7+/v7t7vFw8A7GNsxX5ZF9mLpp90zb7fc0sMp+c0XPrJDNVJ9+cqIjy+eKxg7w/ovE8v8szo+C8t74Q0Vjj6Rsg4WfBpfxY9PXvvauf/5P1l392+8SLO3WhqoixrUxkOmdiCtmtwpGBjmyMRA932wYRtd6AUB/uZmZqHs5cIuXuVGTaiZhYVBuJMJGahrb3Xz1sqWSkTZ3jv337n//Lt3/3xzftVre61a1udaujbgL0rW51q1vd6qPrD3/nf9iKylVbuzu3HJu+ODVrvS14PGaVyIx0TqcMKvwhAbOYnlkhYipyjHqqMG9RVLQ9aoUaNWvFJ+LGbMTKJMty7uc7UhFpxPbVP/jTz3/pz7/23fffe9x26ZlZJKc5lYlJVdrSf/7Tn/7Vf/yr27Y9Xh5P53NvCxGPMVprxAQPZ1ONgEmKm1klresKjaCZZUamL82aiVT2bqaE+X2RVs2YWVUjK4sCafFMOx2S4SGCt65q5ohl5rquDw8Pr169gqUL1OJ9N//dyBs/9tNVM7poGqCLEmBrhu95DtYyUWSy+zHxTe4cUUSaojrH5ysBtTww0dPOiSdtImImE4MeXZMn8ASJ5mklg06qGdO3Sx5jGxg/z8zKjXmGhn1oNHmiDGKXAOcXYTk0s6HOzFD/MUuOXes+iEijng08zyd/uPMgmKpoZBCRqY0RqgIEaoTDOK6m4QFkim6qZkRgw7h7brpdRNdt9TEyCXbXsTkzb9tAohigHGA1HHvjGEKHtsk7C2XXPQWj+pkBXgYkUY9gojmzT0RUkZlU2xhZGREAjOAKoarYs7xkZ0RETP/gug5InFB+0RfhHTIjwhE5BTudnYOsTeGY23HSMFZONaiKiURlztXLZJtEBDGNPZKOmYFCh5gkxLulkYEsyJ1po/t4Qe3EA6QOHjZqmK9FRGRgE6Ds4RwAdQGXIa7BMQa+DpgM2h7MiOPiGV1JVFTrtlVBaz304ulMxzu6P3rkuq47uhw0BlrXNSOJaWxO/ATKaNay8jBQi2jt/ABsbCZ2fjCS9BCXJwLyb2Qelv/r9RqR1owINJiATp07hx2tNSauysoKMFu67gRhAlWmqeH4DXdR3dbt2EvHkARcqNAozWwK9AxSs8C/rKIROdVAntji41ydmzBPkDKo/xFgSoC47e69dVWNijE8IsMTLYp5gGoeov0UQvroE6SCiFydmXf8RZm1Ihrb+JEWgu78+mPx3YYLc8ZkK/E2sIBg7WoeRHO3MLPamD+e9bRS4VJkjCYgAhTNM5/tk6l3z7UL57PNbpyPbeBSaL1l5HYdaH2F54QDTWbShKioCB2MFBVVy0j0OSK8KrF6MPHj4wU+XGIBkGHbNmwLzMXHSRUR4VER6M+omQ/fxgamM1ZIwYLPnEVjDB4+xlCV4wWJqHaH/gRfPLtk8D1P8zcIcCAaPogIpwQTxY9Ks1U5Wc+QxnfxGS2PCaipqhwA7tO0OhNlZAb80ALF/hntah6LcAfh+rQsd+ezZwI/guEMz8hMEa5iMOvrmIbBdh2pvFDAeXb+JhUdd73nb7lzn+tHNvOg2exfsKaq0jKvwpFZGVVBlAf2pKqCuIjefdj+7Xfe+9RPvP7x1+5e+8mPazrFZtYpkW6Kj1rooVsC6ywmADSJSBCxzaGfyiLTiRiCV33vZs3xAaLiynlRuTcWUVmJOGU9X05+UxVudatb3epWf0vdbhW3utWtbnWrj64U7l7jpKdTP7e0Zu21N1o/iZj7FLyuD69ibJzOFfg/ZeJxv/W2LIuaIaGKhM2kN6OMiLEosTU7NT0v3E6kC0kjEhpErCTIEeLLxT//x1/+7O9/4bs/XMOLmYTmTHIFvEzFxK0vb7z5xqd/4Rc+/elPf+ELX7hcLp/61M8Ii0dcHi8QMs7nO2Hmouv1mhHCfH9/zySvHh6gy1qzdPcxelczfv21F9s23Ed6mLal94MGu3lEErNGFkkBQZBZQHJGpuzgSCbKiFevXn7wwQcPDw8fHsilv6v6/FFVsFwVzNEsJOXgtk6qI9Sc2mP3aPfB4ccRuiXCgWSwmIlt1trBrQaPoma0Wi29V9K6Xg8lkSeBZJjZ3d15jAEtVq2BMf0j2ta6rZWJKftdyManAsOBDzgDMvQiQkRbOxQxpWlDwzS0wtLLHDtodNptgXCtmhbp1jreCHmSOdPwsqaWJ601PO57OBHNw/fc0rbTYx8fr6Jqqh4B5CikMcUgtgjvr3+40KuiaHYvMg5+CL169cAg2u5c1KpyDzRagBfPKiZOKoStwfuM1/EIaKI8o+GiMoX5YFOY2XAPD4RzYtgctBz36enDfrDW+tL7slwuq/tGVBXJxK03zASACxoxxR0Whszel0Um2dmBO4BQa2bgrTYzU2PVdV0hGZ9O59ZbeIwxIrwvC4IjDzb0vLTmoLoO0KXV8Na5C/1jbHzs1ayIALMVqYaQ2LCBWBY8I4uYZekLUUU6pOre+7ZtGWlm0Pdxbi/Lcnm8uDuLEDmDhC4MPAV6LVWPkONxTT3WI4zMsvN8AEmIHbYb/lhFWUEzWTXny7LOv84AURk+wmM2gWQOf8zBfNnjCqswh5GVUcRCOu38lRHIWzPk8o1N1Fj45cuXcz3aJfunP8hkz85rTfX5abb07p5UJTr9orkzduANr5xNoKTsvZnadV2pioVph06s27brp8QkaTncr+u6LIsIowMkzOfzHTFHeMQoqknwZz5409u2oeHRW2cWuG73BpuIsMrMS0S64+4cD6oyM20W7hGZkWYK8/LsX+xduslIGWPK+c9KJ1NImKmyInPGkOJfAaIyG8MzU8APQXJARmbenc8iGu7Yb2DjYNFj4szAKm6mRyAB0PAQoJkJtxtrDYvk7AGwJBWLmOlwr0xVQzag7ssvEWVk7J7o1pq7b2Ns23awaObNhWXCryIiorUGbjn6bWNsE7JRBziChVlFtuGRAQx6FTlaLFiyqmpvNoyMqmcQIK4Mr4zKQieMprV/F6CzWm+iUiMC8yYZGKJhglhKNH3QH2U6rnIf27aOcfrY669HxMPDgzYDcOa6re6uKj8qQO9tDHxmKPjo3OA1d5EdP5LPM355X6jrwx9jZyPNXwhY542aWEakb1vNJmxNAZsn0PphUL4f3/3h9a2fldfe/BnLVX3tWgg+VhE1hMEOtAfmXZ6kstxjXRdhPvUFoB73ACgcCKuqJJoxobhTYCZJmFXVq5beivTlul2iPn49DZPPvP0vfvvt//7Hd/WtbnWrW93qVqibAH2rW93qVrf6iPq93/uforKMmrb7RckfPC5JuV0vROKBx8Ya64WqTETNui1Ls6ZTSauMzIABSVkVcfa9UTB76dLYmE2ZmMZK60ZiREJJeOQUse+98+6ffOUbX/j8H33329/l/cmLioqyoqhquolF33zzjd/8z37z7u7uy1/+8jvvvHO9XItqWweel+b4+dgoi4kwyNzMNh8Z+fD4AFrrZb3AMeWFzz+rMjfPy3XN/bmXWKNoRECHxoh97nPvEFjBt6TK6+X6/g/fe3x4rCyieLaP//7V5x8vPKyT72zHvWimuhXBfqmqolAxNKDSMRijVQcwdR//jSyiymImZcnciJDiSEU5Yq2JqqTyePnwQDupWUYw0OBToHA408Ek8VhrajKFeWpLzXIcPmburSEG0MOJxjoUiuoR7zbGYBFTATmiDtvzEwL0YJtyZm6+EpEINw+owzwh0LxFUmUgrY4osqaMRpPQCvhAZqioKEeRD1/HMFFirkz3zEpNESkYGNHkqII91SOiqHoBWRC9NUiW2/UCeVRVmHjdpt+Tmdl53WD6LsCLRRU+5NwSQBJmHcM3oqV3YSaS4YOJiRVycCapiKps7tdti4jeupkiLs9H0K7WeGzXdSt6Ba3ZEERZ5OC6crl7Ecne15inNTPICBsoydBcNicmU93Wbds2M+utL70/Xh7D3axtHsLi8J4LP163w1cLREn45AbwhKpDBHuU6aucso6qUFFe1/0AZe9dRbfN1bQpXa5bZFQm2B05hX7e2qhKDycmZlk3x1mzOUbto4j4uvKrxwOJW8mzWZFRlb01EckqWE3bfkCBeaGJQ2EiyIicoA9HRo6qafvFfD3S2LaBtsecuhgbDP5FRVLC0JkrM6uZJeW6rq01FdkZ0MXIwctA5yQyMYkSzPAtMyWy7J7eCIwOuDipYh0TUI7FcN0QL1tUI3xcorKEpRGB4k2MEDfZrrMjRUSAEoOHnlXCsmMKpha8r1ZEJAyICvM6tkNwJCJ/fJgLWkU976gx782wuexctpWK9wbZ/E4RYZr8DfSTfBppi5ljOLnD0L2tmyYuPyikuQuGbB7gDsseYnnUVkG5icnOzMma9lhQmEJcVJ1pxgPgpqOiEaDQDKKxbRvI+IdEua4DJ2RWEtEA8yErI0TBNKfaswhFpMdOY58LFQPtvQ6Zp4QnERVxRo4oHi4slenupsIi123Du+fsrj0VsxKhZ1NUNBC9qApl9LoNRmdEODMjQ0W1tbYspDa2sY0VQwv7sdOsAERotkuZj70NP70QJ0tJqgqal9ifcNZnJDqUJMTFnI6ZpNkqLtjV0R7LZwLvIf8WVV0vFyJWM1MVZixQrfURIzNZGqP/U7sHX5iKxhjQZEGaOlRpItpPRZxr8nSe7qChH6nnX5wmbfjHhc30/v7+lXv6bqcGEX9eCeREa9HXvv2DN17c/+LPv/WJF3Y6seaqxkKt9t6DlgpjBAHXy0SfI1P0WMAzExGXeDN8OavCA3ER87xiVtPI2sYQPb/w8b33PthCyRbaCUi3utWtbnWrW31k3QToW93qVre61UeUsq5Ei9Zd1xiPNa6cW1KqFLNQJhUpky2mKmZNmFTYRJgJnNjkOjyzxOwRHs4ZHEGVbCKsTJm+ZQRnshoS6n0L36KSv/6Vr/7r//WzX/2zr73/3isiJeIn7ynR8Rj54v78qU/91K/+6j96//33v/nNb37w/geZac2u162yYG6NiLENmvGDTEQewdsWEdvYRERT54x5FbER0+GWrayIYA44vzJTrLJoGyMiGYa3He8AP5O7E1WVbtf11atXj4+PePdnvqd/F+ozTyb0FH2m3ox9drzp3HUJeAkXcRVVgDXMu4QOeiVhxFgE/3T4tCaxEu8IyLWIFlfGrn0IQy8Ym6tqEYEYy7v5EQwQPE/vdt3dq8jgmewSOaAL+xvhe2BuxT6fOktVRHIWVaGvsWfv1ZHHJSpEnFVmLaugDFYSwrSgU8GrqElZSSCMT6D2E26bYQsnypz6pxm7+/ABAY5U1QwqDO+pVhMHzADEwtYK7zmL1tSzateNEPzHAj8s4sWIJk2gqiJTZHqdPSKdEHvn5FzCe16V7PyU+Qcq4LxBoqjENVpZxPsugGhFRMKalQB3qIqp4ohMvYILx2pagIkyEjSL2nPPZuwlq6dXTuEQ2VxFhFkBsiYiGRU1IlOVhBUWbGYmZc4Kx4g9Z4TQdJQzF1EeXRVowaZKTDAMVtWePjdJuyoakkTEivVkVzIh/lYV0O3C8JMyCzpJuI4qE9sIzzOrSHFAb4/kLiJKVfBimxk0ViJWMTXQ8isihBFSqDB1qwigJUCvEJM1w/A75HsiSD+FQ/yko7FoSRWw3VmlwFwQTRI9rrWdhFvEzAfypYuaYkF77tEsFhIyVRJweIqZ1UzA6NiGiML6GpkZCT0ax7lqtgcmKSJ3dMnuoqbJ0yCa8ZtVdcwK6I7ZmXj6bVuBEBGS2kcKdtPzxIgXF4IoM5PnbAEXFrh6+uZ5rHnK1zPOcaeSMB/rHrYXiz+ZYnKCcj/nZ9ysBxnLh8XEzAwPIy2p3TpNSfPWkEkZER6qmlU+nEWMTFiPy7qKIrIm42iuBhFRRKAoMFAeRTld2ZkUTGh3OeaCqOa2HIs9w3D/JNAnMc5EqoqqambQI4uICzc7mmSJyaGhqerOpSsBVwFoIyJp59hUpmfqtOAXY6PdAaMKD1FCR+6YIcEqBZq44PQjqOfzMwCCIVMEZuD78c8qMlsUs31i2PAnLZgpCfl5ggYpbiDPb8UOEMfLl6fTCWMiRSTitSM05lny7PeOnN1pJmLwmg6ruIjk3rHdl6B558eOL0AtPsqRfXzsjKhKFmaS1nrvvTLcB0Aitd+EcEg3onfev/z599776rf/annrE6+9caLhRMlCQixYuEmZS4Vxv6hInrpz430bDyc2bnZoJMwmTjdMD8RcFVlNM9OUhav383Xb3nl1oYeHV/2Nt99+++233/7xrbvVrW51q1vdim4C9K1udatb3erH63Of+52MYamtU7hfHt/tkialzKel996mtVnoxd259S6qY1vX6/XyeNmu13Dv0GBETPDcXtfHyxib0ORCmok1M7XreokYLGxmIlpZ7jm2vDxsX/7Sn/3u7/zet38QIzgRqMcJ497z57dPfuIn3/oHP/fJT7z53nvvff+d7798+VJVz3dn9xngVgfSQUSn6DPFRzwrQsqc0IBMY+STIZ0+g/Hwya03sopMhPURyz6WO5+lj9nb3hscmi9fvnzvhz8cY3x4BPjfjfd5epam4FhT5p3/NHXaCbqlqlIWtZ2qSWQQmvcDV2ArZJ2X3jB47k5ZGNE9aNd4ecxZV1VKOjPxlJAiohCcxUREIqaisIVWFeQiNTWdXlQ88cOBBdgGC9+dzvjXwwC7iOwYU5jkGL5X3iegZzSmHKoBFBlureF1TssiqmDQRgRstrslUZi5qcHOGe5VpYbheqhCVVVgFhMwx0R3d8sY4+HhsarMbDktvfWq+uCDl8xkprRHQCIBrCqbtdZbM4OYDutfZZ1eewEshjAJcWQjYnkCNAsYu6K8LMuyLB4Tpns+n4no8dH70kUEXRAR6UtXlmYNx0j2lMmxDaAw5ltXLa1xF1UN94hYTidmDvdt21j4fD5FZmWaGfMThCQzsSvcg2SqjZm1BL5Tqgp4ClW5wwkkigPx4v5eiAFPCLiMiYhYWVjY1GhOyrv1pqqXy0XNzqfz8AHFink2GzKzqMBjyZYZQUzNmpkd0/FF1dsiIma6bdsYY4yx60dTmm2tVeW2bVDs0CRQldxz/3CNZ2VrvZlV1bqu27a11qa783zGSTh8jDGW1s1sWZaqch/X62pmZiYq1+tl29YX9/etNxYd2wBjBAfk1OfluI3NnW3K6AbCtYdDUheRMUYR2Z3Ok0SVqpC+CCncd9o71rreW2tNWR8eHnLa7bWI3L1Uibl19O0yW86L1KyqLo+X1lpfenggz/B0OjHzuo7zcuLdwco78mW9riLEyNETJSLwdkT0/v6eiK7X6xiDmE7LCeeSMEL5+FVVuPdlmYozSC+C20ACKEFELFJPqA2GvF5U4YFWB87GqgQh5zpWUVGV3tSDMnOCcou2dWXm02nZtkFZre+nH4cwqwCGTqpqUD+fVRSRlE5uulQJWlzEpCI4P8ODCn2B2TNhKhWlRh0BpxE6G34UmVlpe6bovGx21Em1wjeoaDIXQvCIAfFQVWjUSaS6NyH4aQE7mhFJ1ZoJ8wQAFbEZbiMY08g44gplxHB3ZjVrp2Uhokh0dklEln7atnXdVujVylyZ27aBfkNFhX4dlYPfXFVFIqxcEZFZ1ppQIZKYSYzJGWM6YGjkbCZw1fTRK8jw4YNZdM8dPW5MJUVc6VyllEn1fAJp3ruIKsI/+OCDyPz4668D9EREaKIQ/OZ7v/P5T7oHtHJVftZAnR1untMVoGPXtJ8zq/61j9477YbQl+IZOGun8z0Tv3r5AZEQ5fPfJTBUdQ36yx+++vyffPXN104//ROvEUmGR+TSGpoyGMbats2sTAWWecrqvR+pg5kp+20d/bVCS4zI1JKKa2KF8IpK3DSpqlTvlkVeXUPtm+3f/wn69l+3gbe61a1udatb3QToW93qVre61YfqM5/5zOPD9e7+JC3Od2eOa7OPL2bdxIRVSbmEksspvXz1WJl5vV7dXYqaqTD5NoAvSNgbs7Sdxc4eE3uqzVrvbelWWeSVTvD2FC/SHx/9c3/0f37+S9/6zg/8YaMoxiNp0WHoI5X5HP8r//BXfumXfvE73/nOwXTQggAAIABJREFUD77/fSa6v7tnZiFlKNVZ7iMyQXZUUeYW4WMMzJSrtkNUjXBmQADMuoEi2omykoqsWWaSO7TN45mTdlwHz3iljMhtG69evXr16tX1ej3wkX/nquPhdrr7BLIBT9ssC7EwwefNux96ciV2LzPhFXbjIlyuYao7yLUgXEIQNcHuUYAFTLX1bmbuA+a4qYkAvjld1TPiiYj0tRdiGpnX6/V0Ove2RALXmcjIamYiSkwREe5Z1VufhtZwVTudT+7uwyMcWiAzR8QYmzC01Pn8735Ws9ampOvDp+ELxw+WuqzI6K2Lyp7Ul/B2VRW+zsyTy8C0baOylmWBg3UMwDSl2ZMJlJlO5yUizqdTZYpq7x2a7Iv7Mz6eO2xxIkxZObYB8bB2RyoEizFG71M+VhHdmxwoVV2WZV3X4UMw+X744XbD3d35rCoi7B44R/Be59Pp4eEhM+/vXxBVRIxtM2vn02mbwNkfaVhM5zS2muipreLuZtZ7I9BpPcymAA2Cq6iExxgBmZ6Z13UNdzU4dOdWMzNlUdX5tEBQ7r0TU1X58KqCGZ2YwqdydHc+mZq15j5mdpxMhyd2RbNWVdA0m9lyOgPPUofDeV6u0e0Oe34iC8DfoYKOnFmRTug9kMD1XFXhsGYTZtKJKCLvzkvtwYkw8MLgvzc/ZvcrMjAsITLP4Y9/7DX0NQCZtRcvmDkyaAdY4xInusdkf8w4T8Fhhygc4RGpIn1Z1nV94rcwb9uoKlWhmktBuMfOBFeRU29E1FpDry0isQ7s8iC81eU+EEP2+muv4RtpoUO4r6Lzcmqt68yrBEKHqyrOZ4J7V2Y76P7ujLMWu2vpPWLmRgo87THP6fb6xzKng5hm1msmUkPNem/bNmYDSUSYwW+uot47MwUgN8Aiw6LORESvvbirKmZSNSxEc4nIvDt1UTHVbQwqWk6nysTLqpqZIWeShXEeH31Q4KGyag5zUGEZnKCYjGNFzpr/QdJl5srKMui5vWHugeu4z+2FYFXY6rF6Aw2Dc8A9hAmSN44+FUVlZOLaBP4bbIopYWd5uId309a6qsTwg7HAzICuR/R5AzEbPty9SJq13jsRZWY3nR9JtZmcloafzfiQ2ju7n0DQ5KTYy6RyV5kw89KXIsJlQgQAiMHOzsfn3ld7YhKWrMpKH07TxV3HEAkhMDY83DHI4RtQyvnhuypTUUZs1/WVvrp/8YJFrtcr7paOeEM44auK6MgIfd7zOG7xT6kDe3oqvojPvO+A/X3nnoHLPiNmUO3eTBZscWuW0dV6hu/NA2JmsDiKaBT94HH9yp+/88b9vx0PLz95p52H5qaQ0CHVMwvTRHBUURYlibCatdaPXqKIzI7OZFYRM5sadv5xl8GxxG5JW65B1+HF9Uv0fz3kT/4Nv8Hc6la3utWt/n9eNwH6Vre61a1u9aF6443TX73z8pdetH66X5pIW0xat2aqJpWxVQ7loMia8TijMtZ1jSLrS7NmqmsQFZKXGjELZz/didg2Bgkj+6i1Zs1YmTgoISWUSPO0Vx+8/4df+uYf/+l33n2kjTjp6ZHx6Zmc+e7u/BNv/sRbb/3cax978cUvfeUHP3jXxzBrmbVeV+ga4bGOLTNPp1OoCktrFhHbtrkHZqurrLJ4+moDjifi+YQPpGMRpXtGuo/dQ/ykKuPpjWgKSe7j8vj4wfvvP14eh4+/v4PDO4JCptlZPxRwxAJmAfPugMYXp4fzkDaYQXkWFsg67qEGdZ6zoioBImCijBTm1rqKZIaq9ilAK566Z0xWBD3LM4wI2AmXZRGzyGCqu7u7ZTm5jzFGRKgorKC0Z5fhNZe+QCiBN3M5ncYYbl6V4GMQHtdzOSzf2DtZ2VrrvcPZ6sOtGXyXu/g4sbCHHH8IB2OM8FhOy5HHiMO6dM+s07KoalFtmzKCFomLyt2pSkR671nRTKuSReAZJ2LVM47Ztm1QrqEHDXeIC+5DVZF2GBFj02U5wdNq0ykcewRWqtr5fG5Nw0O7DXcfY3Z01NAhAF6DmSBfMvNqq6nene/Af3hxf1eZSALsrZ1Op+4O6f/YbIT1RaaqtNa2bVTFVGDDL5ds3e7OJ6io2zbMZHJRMrJKVd1CZZoxRUQYzmmkltEeI9nGulZVszZcM2tZOjSOsQ0gUFozEYGMB5EXx86V8RWZvIKpTTWzzDQTYWmtnc5nDDrkTJLbk8fWNFNrrffFfYzhRAmUhpru/n2vSlWF0IQT1T3CHb5yAGdSs/aOjogg6bCqwPkFQAMqLY6I7ezpbduWpfelb+s6xnD38/kkKj4m5nvbttqDPSHXXq8b5H7dr2h3x2QAziJTOeI9Gdj0feGAtjUl0QhhMZFT7xCSYVHHxxNVD98XCo2I6/WKH1+WBZ5WHFmzedZxl94WVd1Mj7bccRntLPoiqGl71ijv2ARcltiisQXgPHY+UdE6z2o+nU5Iuquq3pf7+7vr9QrvPD7MDCEkQgsnIsbmRbQsyzF2gM8MP/ihG/JuVsUUjgiNYVXUe5undKSaNmu9Se7ceZGDKXxs7KQWuAc8pFTk7rjGYcd2B7gJdlfgeArrJBGZ7byX2Zc6FnG6XlfIzTDSHjGbWE8ikHyb2zZ2EZOyKiptTic4WgjoKlGxu0eou5pZM12WZcgW7gDoY5vg+scnYdWeNiEhB3RChZodq6Vpq1KsxfCnEz3tJFXDXEsjKyL4u7Ea4DP33oioSueSlznHNWqnWOwrPtRRJi6mpIrmmVQ5QTrEhGU8I9TJlSp4qwiRyqQZHnGI/NM0Pcb2+Ej39/cqUui0EcUTARwRoVxVLGLajpOnqgCcedYO3LvE05FNxy8M9aMu7PnuO2HmSdqurODMLBUhYhGd+Qizu/HUonCiV6uP9dUXv/pt2R7/g5//6Y+1sHgUCqIqUHFU2rPJFS7BLYyZVVRwy/AQ9KQzjoEb3ok6OMaZGRm0y9qUVNoH6SZcvZkvr9cHn/mv/8Vv/6tbFOGtbnWrW93qI+omQN/qVre61a2e6vd///evl3ff+IVz78trL84vTqJkks45PU2RnjFGbDXW9FUqw8e2XrdtI+KefL7rp9P5vNyrdeudCuF0xac7tnYG15WZKymCwmMMplQliuBi68tf/cW7X/jjL3/uD778p1//3kqUxEn85Fnan7oy65Of/Onf+ue/eXd3961vfutLX/ziug1VU7ExxvV6NbMqGmNEZjGZKZIMW2vMFJER4DxKZhJz7x3PgaIQ8SZE4uHhYWf1TuBkuhOVquwSmOyqwdQ5xxiXy+PLDz6ANvT3UkhpwgM47dZUqErwQeNvJjptZU8CtLDO0drYSakEiSAc5izmJxvpk4GrpomPmMFPgLwy5WNV/Ble3aYWmROLIaICabu2MYyoqFQ1AbJ8BrvEn7dtQ/oczFYeLrXraxHrB+8fezgy/OpENIPpIjKzmFSUhTmm+jOGV1VrjZmJCU7jyKBiUKKhP8x9EgkfZSWIuDUpE8LuzsSmkpnb2LB10N/HGD5GhOPp3MMhcokwUNgQUArP8HQANOD8YyL4CxO6GHGt64ZIKKJS1YisjJQps+KkIqrr9RG7YrsMuEMZlmof2J4xRqYxC2IPBbCLKlwRqnp5fMR+r6p127YxTDUz13WFstZaA7i1qohaaxYxxpjpUpk5fKtKqhQRD9/Wbf7gFOzqGC8YvtEBwFGFfy4z13UT4azMcCYiUhHOjIeHVyIQPdH7qYhBRJEBFSUy2IkZu2UKQPtpriJ8XQdO4KSI9OGIxCxmiOoCo32k58jIcN8OhQyfLdYAEQiE7G3bmIRZKovo/2Xv7XotyY4rsRUROzPPubequ5rd1JDdJEe0RyJnhBE98uvY0LwY8A+QHv1oAwPYwAD+AfoBBgawAQP2ox/lJ7/IkAcwRx5LgoayZUrikBqSTXbzq9kfVV11P87J3Dsi/BB7Z+a591Z1sdkiRXYGGl3n5sncub/z5IoVK6BmWgpV7rMGdpZLCVZ4l1LXdTlDTUsuTcibGvzqzKyaHK5apjHnPHZjV7XI3R3OxPF/NLmMujqBlPpSInRDhmEgouvrQ8wWANM0HQ6HaKO7Hw4HVY25Gt+axYqAWRBmjUT6YVDVq8tLr9IxOzPL4xg0dgrqehMfcPdxHC1oksR1d41oBrjZMao980+bT8zNdJqmlLpAGIPp33DSEuzMcRyjDiAENbjrOjMX1cDbu65TpeA4Bzo/jpNZRZ/jdn3fp9SJcJtyHRN3fVdKZiYzTykNQ1+KzhAbgFALaQhgzJYqYp6S9JwiUyIT7Xa9malaVRZvmksa16Lm3zPTaL0DzOj7vusShai9MzOlLplqKRrPka7rouSiU5swAXd6gIZmNgxdCFZY1aNwFk6JA8RmppSYuRuGXexmRFX/18wiF4KZAZS6RMSRTjUl2e/3AdyXksOXFvI4AXYzXDW4v3A3FhGJuAdbuz1aTIuZqYWutKTdbueVCAxryzk6eRgGENWAgHBhElEIPniliDeDuzHqE65u2Q3pJXgolZu5aqRphJkVLcMwMHML5YjkiB+gfKVmCMEQoiRycXExjmPqe3NXUwr3QnP9FrZSipbqUpIkLfNne1i3ZzSaf3rmRq9vGg2kcCo3R42kQIQpxi7cd02eGQ54KGJUrwccpECGv/3+1Vvn/Ze+eO/ePR5815OKEIuEqgnPj37VJKkGi5Q8juMwDPFrx2LP4VQzHtS9J37HWS7FXCMKAewR22CaM5TSQObJ3LR/0p1vStCbbbbZZpvdaRsAvdlmm2222WI2Xe/2nxB/93zfD1ymy0suo1iBomYkokgBFPSj3hhOHVPfd0ZEqevSsEvDvut6ZmLA8wQ4MUFH15FVqesoiY8Hm8aSs+qkZSp5LKoGoXT+11/9m//rj77ygx++dTVmBTtq0vf2H0AkRC+8cP8zn/nMF7/wxTfeePMHP/ihljIMw35/xpJKLsNuF/G8x+NR27tvRKN2XeI55VcwKBEgQuAskf9NUpKApAOeQ60DAATvNSVZ6WpU3DYC56+vr+K+H4nuRrPAdBqsXF8LqaYLjBR55AXGoe9JDayGMMXwOQJuZ3Zrao+VfEZqiioq4kTEFEmQyEpBCEDPb8uzhGlFbTyY1FTDulWYg1FlZlpU+i5AsXG6dr8ORMzdCQU0EqjiyEBKIixFSy2QSVWncQpSakXJ3ac8hRhFvTC4k8QVrWMuJRNR3/XaeNlBqJtRjaDRElNAUQAlEUndOE3xEt71PRHlnENBOCBCACmlUvTq6roUdTdJtRub/EKbonDMeRHnNHlEBJIk3PIr1mvd1f36cDC1kOJlJlUNoDpgIyIqJccYdl0i4klzzSVYKZmsZm4zJa7lIEOmiFW3MULUQ/c8spQtJFWv6sYsWjR4n0rM45QPx9Fm1RQC3NVMLRfVYNQuXpbjMVqOhjSLCCr4rsyaVQEE+ZdAacpuxkQxu1R1HEcWCV3s6KAZnO26LlxKs48ELXq9OlmkMkxDBANAuARQYbLQpSdtZGpms2LHMQQcOCiZNW+lYspl7p6YOH3XI7QyVN1dZDKtXN1AhoraOGXmI3NlQANgIhau0JuDmVOXQgemlMKRANWM4ERM40RNj9hbyk0AwBiE8YCDU5JclIjGaUKICAPmpmpdStwU0s20z4WZgnwNQKbsVS7ImCixyDiqWgQrsPA45aou3XURPXA8HqvGBVdMPPYLEQ0hl5iT0WQ3L6WEc2i1a1nwXpnH8OqVUoIefgMTbGhdKHYQN2FxNwOhOyRQRScBXB9qetUpl3lDJKJcdAW0uQNZ1T38DiUCbSItHpHHCU0nwZuXiGaeeGjp5Dy1VKscPh5pchazRRfF+prdJ9708eMBUrSUogA6c1PT+ljRKVvOBqKiTl7qeBGYeaTq7Qhisi9mIkkkqZaZihszOTbqEoJFkVXPbZ4DnVpEkMyLaBxHNTuOEwEMCsdq8MEdVfvYYypXE1MrqjG305R9nlWm7uqOics45YhNMbhX0DxyciLyKob0U605Vcr23LpYiMQUoC83p2msyobkBsrvaqal7mCo8TTNixCgapXZuYFBn5Cgg957fX3twG63CwV8SckJoSoTEHCDvimJ8JLfdfVUxupZvboT5nSENyBocyfMcTfmJlieEbHHEBEnJkoeItkx4q1ob2LQl6O+d5nfuzi+fP/+y/fu9z4mdhGh+K/tDDBLSYahZ5FSyuE6DUPf9T1X6rdVsLwmDAgkHZE8U7XEvA25c3IYqIAxnE1ml0XHcvy+/MYnyg+w2WabbbbZZrdsA6A322yzzTar9gd/8AdTmbp8wN7ZJzseD4/exXRMbuJEICdH11HXSeo4dSRigBB1zOT17ViSkHToB7dSpqPnI9xF2A6j5cm0yG7gvsPhqkxj1slyGcfD9dUTJ8lKVwf/6le+8sf/5k/ee3RwkIMb6LwA0AR0SV799Kc+95nPvvKJV/7d177+7rvv9cNwfu/+vXv3iUXNtGjf7wAEZU/Vpmliwiz7EHKl7p4SB5R8eXlhVtHVIHb1fU9E52dnQfRbAdDBXKuSryFhETBNKeV4PKpazmVRq/zozB01/Li9M7sD1GiSRNCCRSQ6guhN0iKAW7lmURqAFvY7c6No9TrNgK2SL4VUZWiXNmyX3J1AoRMN+BhAhogIR7JH6UJMQsbjVEoJJJGJA4Aw1YaWekpdEsmlEFES4aAej1PlpAcWAT8cDsS83+0CjrKWgKu2Gq5qItwPQ8nZ1ECV3E0NvajsReaQnkgp7fc7Erk+HENSoJsyAWPOQ9+LyHE8BkidOiulXF9dw10Sn53tp0oi5pS6lFIQxEw1KGw5gv1BKUU+NI8o+IDLAbCwFCHi6+uDm6euy0VBKKWEPnLMSRYxVTM19yQJRGMeQ8cmJl7f9VOeAltXNfNIa+YhAhsdFzrULBxwEaiKCORcHB5iEVSFGtRchSUANUkJgBYlDskLDggkYsPNLcQ9pmlCMI1T5+6qutvtmCue5WY1P6G7qsKdKSiMHPrabp7zxCypSwF/ADiEuDxz35UqeWxmWidhCA0DJFz1ZKc8EVGXuoDsrw8HZu5SN+w0ahvQXhIJqdNxHFvUeeMYMsW8DVybiEvORbXvMxEFUl/Xkru5mVrXdV3fR+bGUBgH0TSNtW4iqDLxzsxdlxoh0tqyiiZweL+ISbOZuSSpXrxg4ncp4PZUokvD4bAkZK0LOQY0hAiOU/RYl4RZACqlhCRxqKdXnN+MhQFysylnM+13u9R3wnx9fQgybGSwDOA49JPMveQIaGDmZCE9dBxTkmEYas5Hc3Ml8uhhwPthMNUpZ2EBwc2KFgBDPwRQ3ZDOJpsMaClBu06hA+Vu6mY67HbMPE1T+GC6LgQcLJBYEQnnRYUwgeoS4BBXcRHWSIdX70YaKQpSinWXc+57FUnjOKopvOpQ5ymLpHDahfNBmCWlJJJLdncWCagOVamAU2fuXvJkVXikxJ7KzEGWr1E3SULXJecS2QxDsFtEJCUCQv0gFleSFHIiGin9rKLE4TObcl2M1WHjKKYAui7FXIxmaqgkh08FLMySJA7G8g+/rAPE7E3QHA4zD3AynDeYFwQMgJu7mjCDAjWuLiK4uzmmXJ8mPnP8QwR/ftBYLIt4iHHTf54FMWYcN0bO3bWYFquCPETwHPhtTG9UHw+CnXzrkbwIcVwfrkG03+/Pzs52u51XB1fVPo4KmMNnfZHGcY7VNJfYPMV1gautZDhOHuhuHJ6/lpuXOSVJSayqddSnNgtB2I0tO0o21SUhRmvDQfHwUL7/zqNPf2L43Ccf9MUSiiQahiH1A4kcx3GaRgZS4q5PwzCY2dBT13VD3w+7HYHMfJyOsUVHytN5I4rJVv00xEkEodhO7JIm7n708PHjg/3a4SuWzr/8e7/9z37vX9/xI2azzTbbbLOPsW0A9GabbbbZZtX2PZ5cTp940dnpyfvv2uGhH68SfJ9S1++Hvk9dotRx10nfkSQjyqqcun63K+M4Ho7Hw0GZyzjRxRMr2UoWMiYw4frySZmOHbN0LIkTeUCexNjvd/fu7ZB2D58cvvHtb3znjXd/9OPDYTJdXhR99X8Q0TDsfvMff+lzn/37b77x/cNh7FLvIDjlrGoR/m/HY2AlIespAKhhG1FI5bxZ5A3jvh9COiCu6vsusnsRUdelvhdmcTct2nepvoVWQnbITYCZLy8vr6+vp2nSUnwF3f7URo19TMEQBAygCkO3eHesGViNLJ0pB6xIvMT5RjNZOHjRswbBKleVw6xyqxewu3L6iMi0xGsxrEobB6ymZjCFe1CuiEBFov4Rcz3mXPU0VEMn1E2JSLrOx3GmoxEgkV8rZ2apatch1jlNIDocjykJgdRNi0b2vzko3t3scSAv7kCXUgoKrVlR9YojVCq0Hw8XlxdoUCAzTzmbey55ylmEl9RqgZsXBaGzRCLTNFUhWkl93zGTueaQ8QUCIQ/oCoSKlRMHyzLghuA25pwjxD4kO7ypoAbYGkhTTEX3QDZd7WBRgrAwT1MGMAxDgLdJxEPY2JRAwjQeR1OVrg9Z5siSt0S7o7ox3D0JpySROC6otZXqzpQSBw0855KkAhRTzhGQ7iF2kZKq5ZyFL1mYuM5et5p8MJKkRVBCw3DqyiQmOlIAbcISwB8I18dR9aBaE5RJSsFhr7gb19SXZiZMSZLW/tOUUil2dThEV+dSgBq+EN0YgFR4jDiJ11iPmlBO1awUM++GvgLoWrzxZNuEOQZYHahleBhmWVhu7Pi6XVTNcprnc8ka0FXzacERKVStbXgN5IqxFs65aNFIi1pysLw5dZ0WDamEQKLVTLWY6dl+X2d1hBpI9UlUmXuzcLZNUw5PzvXhiOMIojxNcd9AD/N4BLGkru97hwef1x2mFjM8JsKUZ+mhKifsPkZYwHEqQYhO1atRHXXFRswDEghjQ+uq54wphJTdXNXMNKuJSC45XAKh5ODuJRe4kzDAK80mV1UWTl1akqCGT6JoCOW3ERrRxBDGXIgoepiYKRc301xIMq+TEHqV2jdVd3CqPh4iioaITA7XoqELlK+O1TuYxNRKzpyEiOCIp0ZsykREUjPRzQz0mPaRlrMKtvDcKAccxzHyu8ZyCP0lK+pMRDTm7CHsIAJqLjl1LZq9MHMKiRizKWvsQlVLJQFEHo4oIiY2a+D0ChVe/u8oaJlpmdkjDCWyQdbVyjVB4uysDQ8rlid/ewZRhaCxmhGBzFqExRCIhU0jYUSbdZWxPE/CZzyOGwatZRoPF0+evPDCC/uzs3EcI1tinJEWXYoqVDK7byOwYnlgr0p298imGaTtW3duGzDqLGuVh1UpbQpPAYV2D9WdDqv2OGBAAR4fjl/79huv3JPPvXLvvjCxQK2okWpiEsbQd8PQheMn6t/3fYiV43AMERuXZMT1WR97a9DT1bymiIQzjEhrFgQhWJ/SJ+6fHY5TJ90n09uXeXh6b2+22WabbfYxtQ2A3myzzTbbDAC++Qd/8B58f486pkRWDpc2HfokQ9fvdruh3w/9EBKiQSgzKuSmZWIkURuPV/lwKOMEFiPO4+imROj7jmA5T+OY4Uh9R12SjqVLNWYZ4MRd35vx8dGPvvo3b3zze2+/f9CxJh4MTpSHwERU9d69+6+++uqrn/ls1/evv/76k4tLA9R8yhkgq6+oFHxDImKukbbUqI4RAB2AoqqVoixBdapXRIb3gKjMLAAyq7K9Sk3fMWL5qYHaOefr66vH7z8aj8eqV4Ab8bY/kdGtz+S+ICr1LR+AB3+0AdDtFXcm/DrAbuRMVtECM7OABNyX0txhRuxgj4BkmBE1UKwRqKtypxlxEKBBbq4VbnOPoGtHiIEwkWtAVAE1Rmx7IJJwJ1AA0E5VzmKmjUWob1A9yRah3no8JK0DcirFzaX1znywdk9o+7oXVfcaVB7SAUmMqmzrzTD2Ok9CFsObpHMAJERMlKF2fYxEdKZuVoqaCBw12j0qGfMxGHDmLg1qaeIhFTEPhKJx5mq0eVAUmTWYZyG8O4PFZqbmII356THhuQR+WhOOgUopgVZUMruNSVKVJWnVC1GIBt/DEtscBu8oWmUQmEgKi1jofQurFEkpBcW5aIiZOtTV3AxqhZQkiXtg8R5S5hWkqtT1OmeJwMyudZkRh2RORRUr/RvsZG5NsLxYIFOhhFFZoDE7AsYljmypRTW4qIGZasx8gNvcLkWDTBnyCTCoOEAWkLe7F61B9KYhLB4cZKaQhbXGGIW6hYqEqXmEj1TNaCOCSPz2dqoaEihaK6Nuc3/EDhZSLjOCT2SkxMwaTESQmWkxwIt5sSobnZJXaDWyL5ofp8LMOWtoJ5kpk1N1kLi7ew4xa2ViYsxzPRa9GzR47k7kMDXPBSGb6wFAq0UKPpA5VKsmMmpMgrs5yAlw00D+i5q7m3oo5VpNztbQZ1TXCFCxQXKYKxtVj4n5lAtHC0Mu3HNL7FncHLnyyb3tlG5G6hqp6kI5RGruWViblFh2bIdTeMjUEY8ENAFidfPY4Qm1CwjNJ0m54aNed9sSl6qBjAmlKAhErIbq8ChGUc1Z1AUAOUf/w4kdDlNlcSK22FDI4BCB0+wlCtEeiIu7myqbxAKPVRbMVgDmVn2UIHjoasGtPnLdqal0UPV0+uynbM+ixdpjqn2iJhiCegd2kLq7k4VsFAFEVuFmnlds4O4Oa2TlAKPJZwR6hl2rqwbtjhTuqPptq3obiblP0abZmj28NMzdSsnX11d930sSSTLlkqcjRyK++oBlkdBpsZC4if/PD2BvYHdoBAHhyyNinD7W527z5puswUBAbCsR/0Jm5OqhfMbesWn4YdxtDoFwQIHrrN9/7/LbP3zvtZfvf+YT+/PkKMddn4eh64cu52ymXV8jVFI6Aku6WnZ0fR9RNfEYrR0bGilVdEvNvDpKmeNXmgiSO/lR0IsBpbyVX+hJf//V1Uc4AAAgAElEQVRf/M7v/sstG+Fmm2222WaLbQD0ZpttttlmAJB39vKRH+00pV1nV4BK192//8L5+b39/pxZEkuSBJ1QjpqPpqPaqONoTDR114+vjmMGxNJgTteX18wy7AaWrqheHQ8iwzB0+/vnu/2u3/XoIlEeQQSSvOumR1dvP3nzT7/6rb/5/tsHwDBrGwIISeP4RJ985Ve+8MV/eP+FFy+vrr71+ncMHkrBJZfcFemSsMy8pFmg1t27rgNBTYs6aRYWJ6iqZUdGKSXUTd1d1XJWYmKmnCuYmPNkpoCzCLMEBWx+czSzi8uLhw8fPnzv3QiZJZGgMH2oAaFbb6oRizx/u/qnRihTfeUlAlNDfwhVHAVe2WG1cFePN8+5fwAQCTXWGJGgyYygxRSLsBZVVZpjxmd1D5bblcb8+u9gibRjFQCSmbIdkJwa06qNRKhB5Qw0T0QwoznFH6ozaMEkANgbZRhEzBISBYCrunkG8ro/iaioQSu1HGAzN1NA0YAMU1exrusANiseQsmJidjUx8OBmEVYUmeq05iJfZV+ykPJl5irwAOzEAeki0BjEVxgh4PBtavc3ZyDpeoEwAzEAqBo5VCbOXNioSlPgff1XZ9SCiWBUhTQyIlHxOqWpzLsBmbOoSDj3ljzAOBkgIdaQQTOq2PK2RtqAuJAEYsZleh+NoW6FSspJRaBobGxmcUldcWUKpHZ4DYLnTYusLSlSrMF1F4ldVPqug6gaRqjlyNfXClFRByec47cgvM0nmdclzoAlZptBmIQO1hSnWC8Zl8DvXReoUSNWIk4TTpZyg1EnomJkiS3bKaoGrWVyc79rLBRnUOMFA4iVyOWLrQmrCG/AAlLq0m7E4FIeLkvkVP10EDVQczC5nBiShULzEWjScUcpq0sJpGpOEFjKB2IWU8zUAjPAQs7m8daq0uZU+V9q5rDpN9HoVo3ZokFxomj2NgE2gprjarr0wHn1kw1cwex0AI6r9cmg31BHD0EY0Ixg4lBLDaDpE2jtl4sCeReNDx2VYCjjjO0WO0WgsVeJwltg6HVQCy7a0wGrzWjNO/DS0tjJwqqbOhsUHiRiCDsbgCBOVTDYy2j4sLEnFqzQU2KoU3M1pEePOjoLqoDF+oTQXCeAWOK9esI3NrARJy66MrwY63kIVoTJcVsbFE1REJYpIndySnmZYCkTbFm3kMWq9I+p0e9ampwYq87DauqA6nrQkoJ1b0dRGawhONlKaPmMVSLgJjoQQR8TgRAhOuqstl53X5DrCYXwKjeyjuezqZlVL24YIe98MILpeTHTy5il6lDw5K6vvK159lCRBRLObykgeG2YW0BSetlPiP30fERp1VKifOZxdzUjD3WDjtZDQToOnYrbm4Bo7eWEkbHoyO+9aP37/VvlP/wMy/t2K6fnA+yH2TYddM0TnkCEL9hAoZW1b7vRMSLEVPdk4WlxQQIV4GpiJsJTZ74fSXSSRIWdMVYvJD3IC6aBTqdKa8fuJttttlmm222AdCbbbbZZpsBX/7yl0c6lAf64m6/Pxv6acJwD9hJ3xP5cTpodjiECWVCGckzkzM7EZdcDtdHB5+fne9258zJnc6HM+5S2u8lJXe7d/8+9cKJO/aSp8urS4/UVGZZ3TlJt/v//uJrf/RHX/n29x49vi6lwQWNDuQGY6pChK995rXf+q3feuedd958882Hjx5FoqTjceq6ruu64iUAi5R6XilOqGpN2lYzwsM8sud1QRMENT2EEFtg9gCNLNDJyJWnZiqSqLKBgrGLwKyvrq6ur68ldUEsdS0fnv38TJtfXFfwcfCu2nv2jNa6B0J6WsCCDiwltC/ikK9OXV1H1ILBEfG5DZz5gAoTcUcVgwCYmBOfQAv1XrewjLvsDow7quxGRNLJ3DuoGtwVJblR/gzBOBhLODr5IvBd82KZFmbeD12cETg1Ee13PYCg9wpT2vUzoTf+bZImVSmCmFwNhL7v4DB3cyOiLnUVdCTMmhjxhm+kgVHVJs5Dz5Hpkci7gN4iAR2AjpnFAYgQkwuBhNNuYCbAO6F5Yc0DkIi7UGiNLGpRgYiUDzYrUQDLTIQ1iAIQkRUF0KfkNUefecs9B0SCLb8pvOoIOeXo0IrOCJtqJSkLm9qUsztKyTFtYi0X1dDoUDVz14U3uHgp8pQBREZFcyeCEYFvQYdRsfV0X80SD6JyBYoXuRKwxMTnKlALmE/j0d0RCA5XZN2b1pARKrKvJXo5BBNiPfgdgN3SyZVL6jYf8dUSJ9RUaFhzPdupbj47b9YrrgJX6+1iTWWtVQAZVU0MVTc39ubpWsq52aHLQCwdGenj1oDfrKIwM2sbg/SE2drOnA/54pZsh2lpUHzRqL3V+1Tme62+B4DZr9mEhlrVo8eYEI31xf95V4vXveHrDy2DgVPrFQou7wfYMo1XJdevGmzczvGFnV3ZtrQ8Bqjekal1Ijc3SmP/r+5XR3qZZXRjQqwa+KzaG98Yw5nM3txMgdFquElcqRHL4QVtL4AW5bVihdfKhbZT/cZDWL8+jDz8ee4zHG9VbF3cFBHa4LMe8wzgrltIseCmcbxm3u92RNR1aZqmmhfUAbKcrTnR6pYYwiZBP6dKvkecDp+bzyIRXjQT/H2enFQjbxQN5Z+7m4jA5Fpc1bXUwAWKfrbm0EPsRub28Mn4+g+evPLSof+V+5+49+LA1ve82/Vdl3Y6OIFZmFM8y4JGDXeVwvFzoXoFY+BABDMvRVMiLSXnnMfRHepGLM4EB7mSoSCp7Cw7SPMODPn93/ud3/29jQS92WabbbZZtQ2A3myzzTbbDDu6ft/PXvEn93bdYCP0mqkwu+pUdMqKktUtqJiF3frEKaWgeRIXEPfDbrc/25+fk8GLDqkjERn6YNGhE+/YyS2PJU+H66ucs2oxM6NUlA8T/uzf/tW/+dOvvvXu5WEyoyreiTXKQBiG4ZVXXvncZz/3yU9+8vXXX3//8eN+6IlIzdwbIbdYC8uuHMCK9lilTwEghjvUNNhkpaiqibR09o3pVkoOnJHqy22lC5k5QCFnqWZmWkqZpny4vlZVYiFVx5wf7Dkg1ee1Gy//tIIQ2yejCrwSkVMVuHVeXUsLaFP/pKUAqkBoxXlugMQEM/JZt4EiAd1zYBJRxYWjR4Hv37jSnxOBvrNwOMyJGcxoehoLxYxARL4qnkBOc8N9hap5ldiuUE9AsgYRlsQBR5qpKoFS37m7qVqT7zjBchwI1QsPhRS4h3irkyQAISnOTDMjErX8BnQSuWlgtA6qGOEc1G1GzD7H1AcSU1UjDIAVh5mWAjixWAlRcmqA3jJ7mIhY5oVS9amFV5A3wQ3CWIDOuecjLSe6LkVYestX5sFkhNyMPG+AZ4VmAuMGhdenLlIrZFwD+a3SRjkUctUa5lyXajhf/HQYK14/nxOL4sascW/qA80WcmUbR2+GRmwmZg02rjVQ1l2nydyJGZKq8nVNDmexUkMNvFjBUmDlIWPWc1/Zyd9B6lzXCnO7mBqFfFFNmMfWAt+/0e5bW8ktqDF6zlBVQQKAjtCK9bl3LdcadoB5oIGK+p0i4Lf1cP30wHKOY94sli3v1oeKxwd2F/erdTlp3RpibY+ZCoquSqw6EHVO+dop+hRree6C67sehbpsq6T+B9hyt1XRS8kxYczrlAnFY+cql7xulNdvnQjO9fImu8N2shycVit9geJvzornCOepD6CTq8yCLdz6sGbSjUmhrpXl7rWGnJIT3Kx53pq7wuNqahTzVmcmEIOJEQ+9eejm4CkCMcgRUSaV/8xO62eQh6MNQDCDp2m6vr6Wrt/vdtM0FY1EpjzjxwDE2RpwbOaz1AlFSc1rWNclk1hNltAU5OfJQvHUjScXCHW5MUf6VhaxUqwUWKH5BtQe23VjJwcp8ORYfvjo8L13Lx/c23/qxQcD531P+30PdA4FEZO0MJ3wIBYtqlaYWEQqdo72wIHDnUBdSplJKB62pgaN5070hzk8d7JLqXtiVorKi3vN0wdPmc0222yzzT42tgHQm2222WYfd/vG//2/Xanu6D2hri8HHN67fPI2k6VOlERBGnGmDosI667vduddv2PpVK0b+OzFXvokfaJOMB7Jj+IMLX49xasZ3Ow68paVnHOepsvLy5wnAu49eOV60u9898df/ctv/fW/e+N6rNLMFbutb3OV43X//v1/+p/8089//vNPHj+Zcj6/d+/lV17uhsHNLy4uSy5qag0lBgDQKiudYwmJJWLWUtVyA1OWCpORSCTso3E8Rn6qeEdNSYrqNOU55L+UMuXpeLwuRUspqtnMmRqfi/gOpOfD2+2C3NeATUUPvPLuQvwUUCPDDLNiQZxRe2guDEtnE9wCM7ujIidaAc8FqVQLslVQvXiRTD0p+aeB680RAHRIMFeS5wxSUosNbzdb+OOVdefuRGCWrCXQgZZgqhT3sb7zMwfyDljJZuqmxMlrOUtjAIdqICOIGPzWseOMzjlmvKbCbSu6HM0A9JrguWpAXSkzTY6JSUKiGwitCLIyOQAWWIYb6M7ffic9H2CoTQYiBDjuDtNMN0FDmv8H5EOrR8teGPPH6DbveGEaetQ2KOp+AgcZTrrJmZ2lltzuFEriNypUKwyAag63m76O5ayb1OybQHmdMjP074Ar6DiNdXVzw43cQXCjovPUumv5r10UJ0eeTa29G6utgGsDjLx6PlbKBXeQdh1+s2IE3OgHDyzQUi3ZFO7zrrK+dFW35lNawZezt2O1BTUw9652ntbhxiIFbi+DG3UJxeQ5UAAh6U8NDY5hXGqy4oCv4NfTStzcpp569xku9xnGXeav15nzXEXdAUHfKHm1K1DdNxpMuwKgK6g684WBJktkN8tfPR+wvvzGSWgI+VO7AHcExczLYaWI0R7sKO1CeMwgc0EDoBvyPo+cV7R2hvpBhURYuA00In1fNHMmX69reLv+LQ6ChQGoKTGb+6P333/pE58Iva9SlEUAJmKEwnvlV0fEiDNzGsKz6Fo0fI1A432H1rlpeLIW9BkgIhE2jZ8o7cx4BDBbQ7QRMRycwtnpNZbC68PFyb06To+Oh9m+++OHn3pw9o9/9dV9V84H7M4TsxF5y9VLcV+RZKqmGikumSt5e9FXcQ/p8CRJtZRSInuHA1ldoxwQg2GU1SdId3V4/ziN15fi9Pv//Ld/93/810+ZMJttttlmm328bAOgN9tss80+7jY5n4uNLl3ii/ffLhdvaxn7PoHJ4U7EzH3XJ+kqPNsNu92epSdOKVXGoh4nTKMkppKRs+bJSraSp+norkGpCXox1BLopRdfpJSoS/3+xYfffetrX/v3P3jr3auxRPwqToEKAA5/cP/+a6+9+mv/4B8Y/Ovf+MajR4+yFunSdHWlahFxz8RqJSAtIgkOUiVZqgUDMnQnuQksmJqIpCRA438WE5au69y8lBIvlpISVdXV+uKoZqol3semaZzGYzA3G1BCt1Gej9j89icHggSN0KOo0bO+gvJucJ/JVuhABTVxGzBa2UIyrDjXByDQs5LrcsQN+hQQ4wN6bPn6JlAY9XB11UZ+XJiYtZonBMuZc+poNMf4YFRmzlrNk9ewDycEGzG486qlQW15JSmwtBMBrXrjqs8+iRtCAj7/jxpqGWAfeUvORjNIDSDA/Jv9Tm5w0rkWVqFTXSrjwZB7mtWhnHGHoCnW7+w2Sbf1XZ0zLfWcc0NsDYCT83xOK2HGSBtgWQHUGwxmrGanWyS7jD4KUd0E04W4ukaWPAD56AvHguPf6LI7jp56WBqUWbmAbbbMvEWvWj2BAVUBhBXsWju/3WdGAm+xSe/yMayqtsL6aZ6vtS9uCBXcLOX2sN1x1q1jBrhr8zC5OhzOOK3SrTnhp4hzdMa8Ey6je4uNfkclljAFrEfijutWi6mis3U9Ey1s2HUx83K9WcRT7AN3cmqbTBROTRZ6abKfnr364wbsPmPjJ3vcChhua2aGgmu0x+JEXFc7tvWZ+WvzHD6pxrJV3nSM3LJn90VssydL6OQRg9ZXc3eZI9QkogmE0CmKdbu62eI6aHFKbRyJ3YRa2tVT90bbhebazAv55AFXp63rHDgVz3OM49gfxxfu3y9nWnJJqSNmiyyyVgWplgfQqjg3tUU2h1CDZ6ypeFewPDS+mLlxopcADF+enjC3LqWYXgR3s2k0NQMTbI6FqoRwhR/Vf/To+nvvPPnxoye4n5jFjjb03HX1pw/cSZhBwsxANJu5MqAjGkY4hZiQicJdRLRwOwcOiLqFoDdCFYU6td4onZ3l9x6WwyTXl5N0z5wwm2222WabfYxsA6A322yzzT7W9tWv/qEd9DLzrifyfH11WY5jPyR0A6WeiJjAwrvdrksdgUDCknphkLsVlq6UfDwcSsmA9YnJQ6CgmKppub4+mGlK3PepH/q+HxIruZ/t92m/493+mOnR4+uv/tW/f/vd92s4J1Yo3EL38ld+5ZXPf/7zL7300vd/8IPvfvc7WQuLEPOUsxYlUJJETGrWGM0AKnwWGtDBH1JVh/vCynQWTpJ0fvM0IyIRkZRY1VRZOCURZmdmkZSSu6uZw810nKZpHPM0AYjg6NW78XPy3X5yuwNC8qXXTg4bTmLw5zOoIWULX25GH+4iiS3XNkh5eUF+jgo3CjBwNwISxz+guAYZnFauwaYMd7gSsYNW+EJr2m1876QswgkmQa2NIOIVZgFHpBEjNw2wdg1xrLqujYg3puJJA/30bD+9Ou5F1LKjrfnbtSxf1xwNkrJ1Fy4t9gb5P8WvgCZYigoi1/JWggt813V+47PPTXCvIGtFmhwIemqc6zUz25qwuQLsWpeti28ADQiwSieve8aJ2wptbjXtXV/cQrebffL5VCUcM9ALn5V85zvV296Asai5MtrSWvORW+mrHW7de7f79wY4Gc3yZZac/rM65yktxOrEZx2IYxFev3gX1i6BdtVNce/WkjXwetdOeDet2G/+cccGc5ukfDIsNx0IPq/iD1OHescPtJN10Jq8lP9BoO36j7UaxrNqNR+nW9227Gy0bLnPrvTtI895ye0T+OSvOzacWqXYFWpYDJrOEAimIIBuyzS1PeLGrHBzGIib4nqocdDaqeVzmMIs93EDfXYAmKMrAi0m0Hg8JkkPXnqJmK8Phy4lEBUNLROSyheul8SviPj9YK4h4VV5yoC7laIBN1eqMVEpxR0iYrbcOgqpSQKY58yrIpEMwLUU0+I1DcXJY9EBAxXzh1fTD967+M4P3+FPv0g0XI/lfCf7QSTEwQERSalLXam+d1NmCQ3o+MnUpy6JsIibA24pfko5FmUeB7xmzgScnAWdgLvu/m54fJgu+/Pk+X/5b/+z/+K/+z8+aOZsttlmm232y28bAL3ZZptt9vG27LQXJqTdXscnuwe/kl56uetFmFmoS8wUCIObqpWS4KRFj1dk5m4GjOPxcHkV4qfeDaZuoDQMkrqu390bziISvx/6fr/r750DpnnMl5cYNaG88foP//Ivvv4Xf/n6u48viZYXzNNaEgO//mu//qUvfendd997660fT9MUIhdFCzNJ38VLrzuEE/eyQj88pUREx+ORmbouEVfN1GmaIp97vA+nToQ53vCERUTu3TsPOY/IyjNNk6qdne/7vnf3cRwPh2v3Mo3HXKaZ1bVSK/2o0ee7Qef15xm7pPoaSwuK8/Ta3AYd6E7gZznHK8es0fye2dKFAHmDCHkX4vYBgHa95DZ0XWGLBvnRHXjzs3vvmX+63aBPoyabmmHiZ7ch5rQvPbF8s8yVmxjqqrGANxVdtPNvy6/g5Pu7a3LnyevjJ3AVnxy1G2c3FYiTWy7VXniIlSmPk8W9mgNOd03u+dwTP8ECHbkDc365m1c74E5uTX7mBKFcn7akbMN6qs5HQpK1NXHW1mg82oC2axk0S86eoKQV2W+E9LlsulXzm8N1q2HR62vM9ynw78mB50Cg7za6c77eKn3tVLmz5OffCZ8H6v2gyJI72M1x+Hlb/XynPfXWwO2n2LPKfFrFnrfCfrqx+Mkkm0nDOOmYp9WHnvJ5LvonNEKTBzmpcP3XWmVmb1qtPN1oxbq4p90G7h75GQAlo8B3ibmmYDS35q+6iT6vq+cnh8nzOF67379/b9jt9rs+Z9USTmzAYUXnrdYaa5qZTS0AaGYKma9gDQMVp845B6AcAvqAB0t9cYTXkQuutc/wdKiNSNfR7oyJj8eDuVbOfd1RarSLAe9dXP7Vt95M6e+bn3N+ctb5kFCmiYEkKdKlElEkzJCWflBEYtQSx09BAYiJUpeImDCLinAphZh3+50ThY6VMCVJIEkMNiU4Olh5zumy2WabbbbZL7ltAPRmm2222cfX/vzP/5XB+NoffOJBJ8nokCgJOQimxU3Z4ORwA0NVx+NxJ+LMZAorbupuqprEzZ2Zuk7QC3GS3Y5TYhZPCQ4P8eeiOI4lj9Pherq6cnBx/tM//fM/+8pfvPPoYlIjZtKFStqAHD8/O//U3/vUa6++NgzDN7/1rbfefkuD+KNlHAFUbK++7M4wWLNSCkCl5JQSs2lWYU5dfQLmnJvqIrtZKYUjgz1L0+7QUgiAqgYaNU2jmk7TdDweDsdjLtksQKhI9PSzG8GV3QmePgOpOQH1Pqi057zd89hPWvKdJ9x5zm0Y/SO0Z4PXP+3tnuke+HB3+dBVuomaPRM5+wnAuhtz8RRc+wBA8WlFfRBC9zwI3t1g5Y0zbnBuT4t9nq6OnnxeQPGDvv5JB/ennJ8fSX0+am/cZmv7oBF4bvD9F9eqR6h9ijyN5GRVU9ktfEXP3nnoxhcOc8t5urq8dKDfDfn6MI4ZLECVUZ5RX3PXmuSAmNRd3U2E3UP62QBa393cc4GpgiAq6698rk37QdOSLpqZB/+YhUWEWVx1UWPBEl5hwJND+c47l699tjx4QHunPUkSkp0IcSepinS5BwDNzNF/kQXW3WFQGJF6gMu5cNOaB0CEPGUQjoddgakrCMyUmHk4n6zT48GoQyER+f1/8Tu/+y//1w89upttttlmm/1y2AZAb7bZZpt9fI21qCTu8OB8n2CTdXAzKzmXMk5eJhOQq3uRoVMr14dr73uThBmANkuS9ud7c2dJ/bBL3cBd712qJKbdHuZ+PD55/zBeHfLlxfH66nC4MsMh23sXxz/64z/7t//v145ZIRJquyfvhOQEeunBg3/yH/2Tl19++cnFxXfe+O7jJ09S1wHuplPJkVC+FAtpQm5CBU2RuUapMnPXmWo5HA/MtNvthEVVj8cxdZJSIuIQdIY5R1odeASiogXVRtBsLlMkU7y6vLy8vJwpSz9vuw0KPwN0oJ8alvr52i905U/s+dDnn4t9EL6LX/xxeJ6u/8i03J+nGAc+UIjmb+fOz2MfumLPLdWz2WY/ud2a35U+TOQ1r18wlm+hz3csjJsYNNzMHj95bMBLQz/lchxHYiFiIWGuKRfV3epvjVMuugsCOK78bABgpvj5UUpxDw1o0aIOF5Eq9x/oM80hW/VXjapFpmERCawbxBUvXm8dDgOuspUn/u5BXzO6vzs7O+8enPVDn7qUOFTIglvd0jmoFtVIkxiEcTQRG3OPfKvxpbm5w/I4uXnOOWuedHI4kSeitDv3dI9MCUDf7fheRv5QI7vZZpttttkvlW0A9GabbbbZx9T+5E9+3y0nLZL6i/felnLJejCdTNXM2UzcCFrKOOWxOz+j1CWGwws5pY5oYBKGpK5Lw447btGccPcyjpaLqcrx2rQcr66uLp7kaeyEhenB+b4/u//GW4/e+P6bP3z7+vGlGmreIWrijo6qobDf7z/1qU/95pd+8+Gjh1//m6+/887b45T7YWBmYkLoJJppURE2S0QwQ8vnA4BVi5mnJNM0EWHKExFNYwbI3XLORMzCzBx5gkyVHMxc38K0REywsEgSSQluU56uri4vLy4Oh4Oquv0t5xt8LruBW90gnP5s67K+9Udf5B2ys3/37UOzzT/Cqza7ac/Vj3eBp3fNQXc/EcC98eXTpu1tPvVzju5Hqmxx0z4wzOAjKO5D2fP5DH4OpX20FfsZ3/G5inrOsu6KF/lwDojn7q47im95MMnhZPAVDZxule43/l17ndwdmvN4PBwO1+dn+77vH19cwd3JcymuZmaVrcxULzAHgwjjOIEWPaIQvI6fOaqmRQOARkJKAqIItJrrEOoqTMzCXt3pCjMCkqTISsCREtDVW8JhAhHY4QVu8O+89faDc3/1C692O04d7ffDICyVUu3mxswh7FH7jKqeCBqn3My8iu24RQIMc7gRhIiJMJUQIvPQMZNup94fMx5N+f2jHvxgTv/9f/2f/zf/w//+vCO62WabbbbZL6NtAPRmm2222cfUksnIx/s+7BJPF+9xudgnlPGgJROo67peuEwH5Im0sGniod/1LB1JIu44/iNhTpSEhBRlzEe4omQ9Hr0UmKWJTYuORyrHZEVYhrTrdztP3dvvPPrzv/jaj955fJiafoavXgwjYRvTa6+99quf/9UXXrj/o7d+9P77j1ISSZK6gZkdUFN2d5EupZRS6jqmkFy0yO3DLKpqZo2o5AMN1LK9A5SkW7+XEshDj4NC+tqUGSF6GG9WzA4bp+P19fXhcJimqcXg/tztmdV47vj/XxD7aDHonw0986lV/hBtWYcJfIg7/nT2s7/jL4x9oD7xz6gef+fsZ9vw59ySN1r235bdDsd5mj1tDH6CCUNPK6gpU9BPIkJyBywNd7c8jZcXFw8evLQb+uvD0dQjd5+7E0HNnEhYljsbHF60EIilyunPMtClaNOXr7rKaCFXoQkW0HMkLzREKg2rALRHbtgQuSaAwOQngVhBknaFG+ythxffu9/9o8++fE9SDyQGEieKBLpwd0opMhly/AZiIoofQk36A4ikkfEbLYjeBDClYJdPWVRTiEgTs3SDu+wLerxQ3io5egkAACAASURBVH30qJSL0Xs+ySKw2WabbbbZx9A2AHqzzTbb7ONo3/nylx/bRTIZdnLe+eV0iXLohv1kaiUL8bDf7XfDk+nAzGfDebc/78/P+7MzkkScQIkoERKIzaxoKWMex6uLq0ewwlaQx46oE7ZMBCS4DEJDEk7dbg/p331y/dff+Na/+j//+L3LmsSnpjtUW2dKYubf+I1/9A+/+IUnT54cx+Ow2336058mFpYEYMrT1fU1EYX0xjAMfd9LSgC06OFwUI0cg4gk8hEf2zEDMPf9fp9S0oiDLUUDqDZLKQkzx2lmasEPqsRGd89lGsfj8XDUUipd6O+IrePcF6nG9ZH5zJ9JfX5h7Gc2gj9tvz/l+p8xIvzs7vp4zK1fbk2Jj8cYbvZztmcnx31uJ+OzMyr6T4I+310OERGVUi6fPD7f73f78/3Qj2POucAtJelSuj5OJwlLmU3VTL1SoUmLAojkE+6uRZk5dWm+pOSipZipJGEKZvGc9RTujpqsQmBODhIO/BhmZm6q87p1EEDe/OmPLsoP3r783lvv8TToGY9XtBP0glAVA5DCsS+CKmAtVD8QN+WxqA2IvSXJIGI3mHrwqMlJKBmsFCU2Ful7kf7syeXV4/ftXjeNZSNBb7bZZpt93G0DoDfbbLPNPo42yvSi3n/M7zPhePnudLzqxCH9cO+FzoxBstt51/XUs3A/DNx1zlyKYprgh1kqwwHVkvPoZmZZdOwEKblpEUIicoe5FzU4m1LRSTImn775xo9ff/Odh0/yscCMnFCzDy7Bp9if7R+89ODVV1+798KL3//+9x8/fjyOo7l3Xd+LmANEXd8xi1Q6M8ZxxDgGicdM4a4lp5S6JF2SCGAt0+juwkxQU5vG0cyqtCKhS5wSdSl1XbLKcDImZmZiVrVc8vHycHV1mfM0y0zD/ScRVb4zor/9U+H3+d35zpNXB2uP0W0cfCZbwe2knCouGfG0RkTE4rNoSehP3t0cmstsr/QtWxIxZuHNm830dmULT26v9KdFzaXVGkS08lMsiGMM1JRJc2sBJ5bleHwVLatEM4845ci/dKu2q+OrD7T0cAx3tNdu90utfKvMMjRucwNXtDKLwpcLF//LfKY/BUCJwvkWvz0qO+fdqoccBoDAs8oDExOzWXGfZxrNrDczIwKRuBf3uHAZoKePzB1k+9Y/c72jZ/ypCtjUzmo4iLk1fOfuziBigJuYqQF8o9x1kD2BvH7gVf6uuXVr3GceYom/V+fPS6XG+9/VF7eOL4vb27xaFkXcgeogkMPjz5BhnW+4bBLedgCaq3Jyr0pdZF4qf6OaNPdGDftY7WZOc/7FdiXNrq15e6nzti0ZOBwna3Np2WnnrEo43W5ofdJ8WewhEctitmwOS6Norp7j1nCsu3fujJs298bzbeYnDVtv23ec2lR91wzbpwGj64lTB51AQYhd6vasqt54gKx2lFrC6VyJWRUyC8/R/Ntr9qRVt06Y94RWG4rpPffG7Y2FcNf+v+pwr48RxJPCb57UeLs3D6+GeNXS5/AnuQF48uR9wD/58icvLi4vLi7VKXVd3w2p79XM3GMzV1VPgupZjycAM5MIa1O3iIfgIrjR9+23BM1VdbT9vz4YYqbFRc7EwlRKKVkyk+VsqgDNyD45yIzcD8f8xo/ef2H/9164t79498fnHR6c75KE7JiFf13VREQ4zSFpbnV5s3Ddd4hZpOuSO1RVpBMWBgPG5JIKAIMTq4PNvaTp6jAWLVY8k9DGgd5ss802+3jbBkBvttlmm33s7Kt/+IdqdjFcdpyECfnQC/VDl/qdBL6jBpHCQkMnXS+7wd1Lng5XRypHskxu7YXS1UrRAhgxeqFExOTMzuQiXN+XnUAJIp5JZbi6Ll//5puvv/nW1egFZPWVEgusQeSEFx88+MIXvvjCiy+O0/T2O+9eXl1Hlnky5VLiZY9ZhCtDp5SSc3F3YmJmN4PBYCEWHfAKCymRuxHMTc295MlX+EEIb4CcGFAneNCMAtEzt+PxeHHx5OrqUkvTavzJ2FV3IW6n790rcuXT3opXb/j1Xftu9BnLq//padRAnwpGExbImepB3PH2fgshPanMXdjjfC3RKQo1Q0XtzXZdd6qvz+6zeuZp+wlOgSg7DA3dXnBFAJF4agEdQMT1T605l056r4HDp923fFhAdvIV4B7GrVet4u0gpxn6b2VWQK/NpwCya+UViBatJGHqTf0WFj+PFAUwuiBujqrFDmqND6w9+gpUUdp6AyZ2kLcxaoOF1QdqSCe1cWT3qBItmN9SLTv5q02cde1XqPqNfr4BjS3IY8WM6uq4gRcvZ3lMmnnU1zedJ1vFdZbxXsGHDdWKDF04BT+rirOv77gqn9Y191uyt23cY/KQQ2udI1faUmabmRRJWL0hjbQ6Pm8Sy4V1+JYaIBDkRX8WRuDq7KCKbAF1pRAA8FLg4nIhAE5ONwMsbnyamx/dyKudgdrWsHjClllx966x3gNpNZeISJbOXYFyqM097ZX5D1qXM5d/533X2O3qfMKCoi5DXeFFb8seNx4ItJwzL6wVMEqndaDTjl1tX1RHYXU63VXCUtCto+u2nyDTMat8WX1065LVwcWZdLfP4CmQ7vqm0U4+rfoN2NpXcurzlsJt0WkDSRkLhrta0afOjXZ4aVtr71yrm4+Y05pUyJuA4/XV0HVDl+xsZ6ZFlUL0uO/NXVXhFB+IwEzMDLiZRY5kIopIq6X0lfPpzsGMW6+b4tVq4mWZMjOz8Ghuaqf97+Qg4DCWN3/85LVP/8qneF9o6KEFkqRjplCUjlA2QIgoshK6eylF1cyNmJujFE7UdZ27aymSIq8HR2Pb7ycAZO7mXvhYqLcyGScxgh//p//yP/6v/uf/5+m9vdlmm2222S+zbQD0ZpttttnHz0TLKNzZS/cfDDgkOkv3Bk6J+8FAqjqWQ87FJiiEczlMueRpOlwfL5+I5wQVdmFmYTCxUBJxgIWHXZ/zNOUsxMwM5iQiLETM/R7dmfMefDb98OE3vvnmd974gQF+QoNCS1nPAD796mv/6W//s6uLy29/+/W3337bQf2wi2DT4zSNYyZC1/WU2CyyybcXOYepE5ETTH3KZcpZSxGWrutSSmaUSyYzwCteyCQsZpZV1UxNVXXK2d37vov3MZF0eXn58OHDR48eXl5cLcLVP73dwRhdv1evT5gRMA/4sL1UMxYs7JRXRwsM1ECfcAsEPZYcHjxoJvGZW+VOKywSdxddb3B6/ATEbPe94/XeqmglASAOJBSYSZdeUQfm2g8cmG9Fn83dWqFrIJJmBDJYpJWV3ED2xjibUTBuUHLFhaIl9aDp6pKFDOvuvlbcdHdYYGPBqXN3YiGw38SipL7Fh9QMEbFQAHDR38yVk77qO/eGS1EjhHpD7ogDgI4Xf3c4TERC+hx1VjgH0OwcV6qZm0VHqWlgrhy0cceMb8Q9zDVSWgEgEuIkTGpFS+2cgFMb4GOVq1tRb4CYmcw0Jlt1BAS8S7PbyWOwguQbVE+AnCrm19CmGe8+AbNOwSNzAkFucDipQtf11gYl8AqMXiHLfqPAul7MjG6CoUyNp0+8zKgGGdlKgbZOk+gu4URERescVVcCM7OZOpwoIYI1YMRMJGbqAEjq+vU20StF2urUYHbzUI1tWwZFejEzNXMHCTMRqWksOWgBQCxQWyAub0uYYI1EH421ZUc66fplSTXwy61O78q6voX01dVEUtu02g3W1m7Iy7yEEXGNcnB3nS+kdv4CE9cq1dk180exvmS1gThAYEbgg0xwqm2bFzdq9EP0SeCANFNWo/QZ+21Ou9O+qYPoJ70Wk4sr0GwhRcXEDHc3NXaAFiR2bmzd5exG1/maar2+/UnbKwLrBBDX/HhUVxnsdFCZ4Lz0KuyU1EzgE3L3sx+MdUHPy9r91gXLc2TtLwMTKPqhJsxz9+bt8AYWn9xmbq/H48DWq7LNgdmFGVU/fcx5e9jHdXma3n//4dnZvZc/8dL14TjmrGpE0qVuGAZVc/M6I8iJOOKo6iQhsLjVHBVORCml2NXb9HauHsSbzW+8b3jFzhvMnhIR911vpWieWvJFW40djtm+/+7x7Yvy6+nsM//Br51hTHZ8cP/+2TAkgquqasmZOYkk9yo+lnMpueSS1cxBfZ+mqRyPU8z5YTeoqZlny6aqpmoWoSrxzAHD0/T/s/cuTbIk2X3feXlEZlbd7nkB8wIHGEgG2pgRWtFoWspMC4lbfQRttOJC3wBfQCutuJB22kArGRfSDpQZBRPJAQUBMJGjeQGcnsH0a6a7b1VlhLufc7T4u0fV7RH04MwG03nM2vreuplZER7uHhn/8z+/Q6c7copoLKn+MZXL/9PMuMUtbnGLW/xax02AvsUtbnGLz1b80R/9kefVtF7W9X5ddH8kb5w9+t72azJ77/vTY+/diUgXKYuVhT1Kr8ShIioioByoJNzOrM07szCfXZZcYl2XxVSF4T7Ggxix0rK+8877f/qn3/nO93/8/s9e/8LRMbMSk6h98Ytf+MpXvva5tz//Vz/8qx/+5V998vo1qkEjIob+iifGK70hOrzxWXCm4RG+1aYqxczKeOAiosjw3pOSWVRtPhYGi5gqlLXRZYjYSnl8fPr5xw9Pj1tr/otayS8R/MaHHX5IPuS2+bI3/sSHJxWPrDxK9d9wQLGIisT4h6EQTr8SeXcihon8ENd4fvSnhONP/eQwmR3yJWU6tGyRl2+EVgDbVymFiSKz98YspZSMIXWIyNR05sM4k4jgjaqKkxCVTIrwWebvLAp5OibFm5jATiGi7o7RGThv1d6ah2emijFkdwDCIREKhwcRmRmuvohkjuPHeB5HiJNVUyIKT/dGmaJKw2GXPHni4LlYMWHG9GMmUY3ICGd8smpvnTIL6OTuOuYhucPdPy40D74NjkhEpbeWmWDRPF//TPcmzGUpvXuEv5wbzwISU46eU+MiBo5QRES8e1KqKIuyKARld58SdihkdIARMkyFoPzHGFY+xMCDK8Bg2sBgFzxqwF2YRSUjmUlVI6YAOo6XIYXGJMYcrHYREdHMiBwCEPEb6wWSypTys5QFOadnmzzRgBzMqX5MmwjHwfTuZmqmVpbeuruPizs8j4yCDHyQh2eGWcH86b1FQHIqIuLesXPFoYiNKzZSCYLERBIxqYqqdXcPx9lhJnt4bw2ro5Sl1XY0MRNmFolR6ZEAzkLMbN5FRc0CalmSiRJR612YMYUiPLozv3FUv7jngdqBlYWFc6wgXKD5aUPFXpYlM3rv0ygpY38YMq58+hccO8i4LDD4CzP17qAHHJtSjnUchwCbmeGuqqIaHphUQ8YemuCYPMySOVT45+KMF6Lky5+jgW2E4zTLUnB9sSHAH0o5mrnNAwv3AE1XBiA4mBkc3t67R2RmKYWZvfeIyKSylIjovamit0HHKJgZdphWKzEXU1FllpwJvBgAqcTW1HtHxqKUwsKU1FpLIjmGbmSPhmCaGabGxODwoNIijwEaEifqCaZaOj6LB+DoUy70PO4UPPfaFFEidncZCcgJmnixcI+EVs4VSWNzeT4c5pmWmb80J3wGq/pYzUMjnVf2OUHIQ15O93DP8Ln2Pv29IpNqbR/9/CMiPp8vrdXtul/3KmJiZqpoNiEiowolD8NyjlFipqTu41IKod3xPJ0kkXE/H2nUfJkWnCObyTzKg3qPzBSmZNZSvLcMFN+M9EQk1cye+cMfv/f5V/aF/+Cbi1mvvu+tiJWlmPGi4spIMR4TIk/jltrDc9wQ03tEBDHJ2Btnxt69R8dPKJFi5BDuog/dpWeTjPVLlfc/+IP/6A/+4J/+DSv9Fre4xS1u8escNwH6Fre4xS0+W3HR7WM/f7l8fFnvte+0PfrTQ0T18BbBIhHeHp+69yDS84VypVyMRDiXMnDLRESiyebCyZIsST1UQu5yIREp55OZ6GAhtuiNa6WMcPvOd773z/74n//wR+9+8rh/6vEOJj7KLGX5nW/+7te+9vWM/OCDD9997z0i6b279wMpuqynJKqteXfK8ZgdU9+CbgIdBupPrVWYTNXKaNVeW3P3wz8oYtAIIA6KyGk9Mct122BKVdOnp+vDw7XVHv4r7T34UizjaXyicQrTCyaoWX5Run44UIfsBbPw4avDM7aqlmIBPSMTMofK6Du010pENroPzQ9kFuKjE+M4QiIiGnLPfBnRUAYgMx0yHE9NnCAK51Ajmfm0rhD1aq0icjqdoLbQaIWkHRLA9LOLqrtTppWCDzFVYvaM59dM6ESEDwGaQKg0ImqtioiItNZExMx67733iFA1Zs3E+yIyRKSUUvdKTOfTuffu4WYl4nliFDOonFCEVcWs0ChYdozGIXPgytAUx5fFRGQK0Ax5He+CpNhqpchlWXCQ0KdYpLcWERCpcb7Dcpapqlas1kpJyzqF0dlhat83Fl6WBRpBBECfoxVnRkCSw1sgIuFEMHnMbK81Ikopk2HyTIl191qrmqkKEWExntaFhSPC0dsTCuDxGzNznIjV1rr7UACJe28iakXdQ5hLKfDVQY2F3o0V3b0f+iYz995lguBRDyEqzG9goLt7752IhFlE1nWdPvHn6czjCAkvUxE1wzlg2uz7vp5WxHa91taWZcnIcG+tQeDDIXlAZqV1XTHC27bhJ8uyqKpDN4pgZohPKkJ8ZLxG6gWDo2allNpa96F649L03iuWsNlpWfe6e3ecIK5m96h7g2S5nlZMqubOwjoatHrvfV1WJtr3qqo2hrS12l6u4swQ5k9p0Dj45n0s3t6JIDICrO/Lsopw652SRO1yPkfEXvc3lcSBjf504oqImPNIQmAlTFW31paZpdiRA8B4DiM5YXPK1ruZmaqHi4hZGWj/oTszVpmquntk0EBzDw8qJR3C6LENmioxYaER0bqeInzb98w01fV0mgbnwSXwSB/LeSxgTCphtlLMrO57d0+ssrnYM3NZlohorWFPa60RkYguy0JM4XG9PrHw+XQGpTcyx3WfXXWXZcnMfd+xd51OJ1GhpG3bMkNEMfpHtojnDDwtK2W21kXQcU77SDsdNyoUmqBhHbFMgT4Oc/QICKYxEydzu3XVwsRtjL9M8z7lISfn8K3nqAPhw0iPfcQ9MkP00zdjRynALLgY9wiR3lp3zwxsDpHxqSPtrXFr7o3CM2JwqN/U03vrn7x+UCtE3Frf9/3x8YnZcMt0zxhqORFTeuDAkTrnyVOOA4+e42Yy7flDpufnzn8875/PryECCYpFxD2QRDMlLcUd2Z3n/gSehC8sf/XTDwq33/s7X+I7ketG7lErX85LUePM7JFC3EVEUFyjKsWIODICNztREY3RRAGZiIyM8IwIT5/fNBjXLYiu3uTpccnyyU418sMv0NuP5dPL/Ba3uMUtbvHZiJsAfYtb3OIWn6H4i7/4w/2T+iXdTmWx7O//279sDx9KfyqLiEowerJTWXRhYyt2uRNbiIV7j+4ZnKwpJqpqRcxIja2olWAiFdEy+/Z53fbsdX98uD68fnr92kSS5dr1X/3J//Yv/+RPP379EMPF/CKYmISF7i/3f//v/4Ovfe1r7773fq29lKUUs1LUVFQjwnuoGoswE5AZlOQReLC0YmrWex+2TWaoP0RpKmrDlt1aPwRoWIOhAR4eo2LGzK+699Zaa9v16s2jOUXA0/ur8UDDLzzhBPgZKApjTBi12aJqz+o03qhDd5bxp2EhPMRhHk5TOTxgU9bOobnASZp5qKtwCyqLqtovCNAw6vKLUFXKhDLCIsUMSt+6rhCG6r5H5rIswyzpPp+xhxvweIGZCXNrDdoJNDhcSspc1jXcuzvOiph7b8y8rmtrDfKfmZnZ9XqFzGpWmCGriZnBaVhrK8Wm806ZBrITYoaZQvxl4nVdDyn2U2ZGXH0zo6SIaL0RkYqeTidmhiaI43F3mN1U1dQiIX88ezYhjkOaHBKqR2/NzFSkDslJ4FGHOnqodkEcU1d+69Vby7KUUvZ93/c9iaCU1v0KO/OyrpR53Tao8MPpHFHMsEDsEE+naqxTLMPpRB4e87Isi4f33uteoboSEWT902IQUsNHUbaKypuWZGImktZaZBy6LaRVEamjUyiaSWbE+Dmc6UTcexu++KKQtCKCKM1KZBzC/ct1Nl7DjNPPiCkq8rPSIwwLJ4QtzPax1pndvfW2LquoZOZSFkw/SIS4lGaWmR7e29DEoecS0RDj3THVHabXCJ6S6jMv4MVfmZkyI6NHvJreSJrmzWdn5XEWxHR4KbG78JEc6lDfWaR7773Bb4vzZeKiBWmYA/kCIyQRASvBb+55OdCx3lorSzGzNrJ6iWHZtq2UIiLJ5D7xIEz3/KqUkkm11pgbwi+m9HBGrXc4f9WsmB1r8HLHSYS359z04OH38N4btiBcmuf6DWbvTkxFB/qg9y6qVqy3zkxq1lsX5vP57OG9e0aoqZlt206UpSxIipgZdulaa0Tcv3pbFF5eAs6o1YodDIJj713RtUC19dZ7V0XW0+/u70WFiFpr4Y7tFzsJJpW/yMnhOnt48/7qc2+pajG7Xq+tNWXGJhATNLysy8vkh5kxcWa+enWPHAmEWhFptbm7FVvKYmaZVPfa/KmsK/6atRLRsp7UDOmi0XNvzIVBKMmDA/zsR04mXtQwnlYWycTxEMvpfJrVNC/eMqYeEzPk/kzqw7CfsEtjlVKKWpE3J0+2lpxqNpN/rqKqGklCHBGqgnT382RLYkoVdVV3896j9windM6gjEmNIc6M3rdtW5b1cn+fxLV1LQsRd3cWjsgjs0UqImKqoyYgx2gpi88kBDPJvKvOpY1vI2PBZ6YHH5VRc/93VV2WMsTfcDVGIifD0Y0gk8c+J8xCTz3f+3j/1z94p/7G5UsrP33y8YNJfeuVcQonZ3hEENkgO3MpZcxe90gSxX6m0749DxrlD2NiCorfeHw14XP6smqTM3/w0etGv/3e5a333/tVfXu6xS1ucYtb/O2KmwB9i1vc4hafoYhN17f2/qGy5fbws+3pI/Yd9fKsWsoqZiLM6ykykyVlcTJmXc8XJrLuYiZmrEPwZEpmFs5I9+b9+jrDPbz1Gr1FbfV63R+v29PT5dXbteePfvLT7/3lT37w4/evteORkpLegFUyfeELX/jm737zN770Gxn543fece/n80lVtBiMlkycya01GJ+XYpQUPjysMAaKys6ZmcUKqvzvLmfCY1o4CakWXRd3771ByXEKVTMrx3Mg9D5lyd63VrftWvere810OmCi/w5PUc9cDXjsmCFRyfTcMZsoi0AXEBEixvPzYcyb7m6V8aAnB4fjpUnwKAN/hnTg9dPEPCqv8cDMtJTlULhMhk8WFjlVYyZ3HxAElmEcxuPtoCVkh/1QBF0imYlVFFoVfFwZCex3MhOFd0eVdUTrLaEreHg4EXGIEfXWIsNzYIuJKckpycNFmBv37vAPOsiVvbkH9Vbcmbn35qEeoSqt9Vor2tn17vBzEZGHezhPazaEFar1MKdxAqcr8FRidFtvzMLE0PG7uxZjHqoxMzfvg3pC5BHdvfeambDEYvbjgkR45mCRZ0Stu0eYGQzCRGRmMhy9nJneezITCYyfHh6UnkG9w6qWGc077WNduffeOzMD/t3dIxxHxjGGTjI4JdwHFEUkM/dWxxCBlpFJzEHZ3VtvESGmLDIIsHC1MmdG987MoqKsEekRSWlWzKy3RsRmNikcPpzdivQJlaW4e3qIqJhIjinuPOjSWhQDyyPnQnBbi6qwyjSJxyBskIhO12QSs4rEM7J2yL2RmQ77vBAN274OSYjAdFZVmqolZNPW23TwUlJi3uKKoHNXD89AFzLBsu3ePQJzyTMlQ1iYBSLj2FeJIglj0huM4r6uq5oxU63Ne4e+JhNGMZD8469jOyUerRNRR8/EyiSsRJnhmWggxqTQlpOZJCnCMTNHAow5I4izWMEg8txBencSERVczSTC/WA9nQjJKhk4ECKOzN4aM6upiiaRCnfvGQmxnsF7Ga1HCTuNdXW3uYfJob+BgwHwRSZNagGB0NK6lVJUdF3W1nu4L+uaGa01U5NpiQUwx1TVDPJ9KWVPYuZlWXBx2UarWzNl4qWUSgnYyNQ9k2HgxpkO0zShAiMiKUNE1mXNRBLHmVhVh9yYmRmcIirOQpyiCk1WVFmYhDllzmRhGrzmYXUnjggRLYWISFkYMwde5kiiLGbQMceNRwRlMXgvfiLrANAXM7Myiy34ENCJSoSVZUG2CduRWXHvmN4AoBSziKit0fMWx0gHttZbq8gLRqAmhmDuhuQaw8A+eUQeGaQqxJxE3TvOaHreo3eHCx6JEpn37t5LJqkqrpA7eBTw5peJyODwAZ3nwbsZHnrY1Vtrve697dEqvcDEY6nv+/749Liez2blcrk0T2K+rGtrvfVOmaKiJjHrFUg0I7w71gMxu4iLH+LtMJSLxMu81MxVDho4dqxhWkdync00M7mPjWqk0X0a2+c1T6KW9MnWf/DOe2+fvvrVL3w505m6ex/pzVEzkhS9uXukufMoQcAVwj1QHIiSkdKG6j2+jxALYFoowsBNpHnzYkYSrVWm/+y///a/+g//Pfpfv////8vTLW5xi1vc4m933AToW9ziFrf4rMS/+Wf/Q3fyj4w0t+tTPvy1cT/fr5e1NHex5XR5FSzELMp7a7X2cOFU4+Xu/vPrsrq7mLAKjfJKp7pT373Vtj3t18fr9SHDKcOzh3sCOeuyFrt/6/MfX/3H7333R+9/8v4njWT0n+cJ10Qw09e//rXf//2/J0Lvf/DeOz/+ETNfLudIT0r35k5weG1Pe+/dTNd1VbXMkAwWMmVK99a8ViIiobptEfHq1Sv33Fu/Xq8icj6fi5kK1VnLP7pmpR71r8P9Grldn16//uT1w8N23cLrG/auTyMi/99iKr80lLPpz4jvWAAAIABJREFUu5xPocyHZCP5wvQ3BJpBFxE8nRJeN9+Jf2FmVcODK+S2qVBTxPDbqqLqP56PSVNVl9NKgEV09whcF3j0TqrM0nrPHE/yIBJAMjuQER0F72aHJ3RZFp6+5kzC0/LxKP08MMw+aQyZeRilVWGrhH2vmBkLvKjdTI/HcyKCpQ7P0BFRay1WWBgP83KAmyN4MHm7aYH6hN6TsK8CI8DzauCS4K3wde77LiIRcd2uZrYuKyyKe92v24aThSgJHkixkhnuDowMEZVSoFQeHmrUZWemiTLRS0M63jjtyABNcGuVaMyEccm2K+8bEcH1HxHX65M3v1xOxNRao+t1DhdlJjzjBzslM3sEc611Z3i3w91927Z1XZm51ppJLGrF9lYjou4DotJnYT7QAZHuve/7jp6fqrrve63VPS6X8+l0enx8FNHL5Q767NPTkwHOPkViECq263VZFkxmqDGDoYFJpcKOZEWKcO/eevNMWEczHMcxfKDLMufV8EofZnOMCQa59w4Pe+/gdaQNTgVScqIirTtRwusds7fY4bbOzAF+6VW1oQEgPhnkDWbetj0zL5czXLHHJ2Da2DT5Yp6o6mFf9cziHhlPj4+11svlDrjzbdsocymrimQGeAtIxeUsbogBmSURsE16a1WHsgpHPNVtMDdwJDwJxSLcaiOm8/kChQ4JseOYmbm2NhqbehBl6x0qFJC6ymJmJhxMzCREvdUxw5lTiJmWomZlpxrhPFkLIsKkpkjShDvwGjxTDCxsMQHTuAIiQqqmmplMtCwLE7XM87q6e69tWQqzuHdlZtGMRGGMz6wgEjDeu7furZsVj97mHAjsPr232rDrYmfLfN41UHOwnk7u3lp191LK3eVurxsU86PUAHth23cRATw6k9wDYmtZCjn16xXJgIzERgEqkRBjvWXm6bQuViLGRgN+fe99v24sXEoRQgUDaD+KZEiqBtqcMi+LDUE/wns/nU7L6XRaCu6DnqRLIXAlKDNThUspp9Np33dMb3fPiLu7u97aw8NDDkQ9l7KUUsy0tVbr2MlUtHunTBEFwQMIF1RvWCnrutba0I0CjOcCPy/2c2aetBAB6zwSDf2YB2aapi8+M3ES62KYWkBaYxdFagGbg4zbR1bE9nR9zK21XzDs8r7XzDydL+t6vru7++iTB2F+dX//+PiUkWJcippp723I6cwRUT2KFbVB6fHhxWZm9tl4wCcfHHeEkYCU55a2x6mN4oNTEWGi6N4jSdUCjW7dE8bucfAcHJv3H7370e9+/St3n/+yLXry66p5smVRFQ6WIArP3Gu/bj2Sw3OvDYZxj57kzAfuJpnH14PIRBWcJ3nkKNoScMOYibI8NrFIIvb/5r/8Tz7/kw/+4D+9kaBvcYtb3OIzFzcB+ha3uMUtPivhwtaSl/Xzb9/7w886nS/lUpSEMtxZLMtKxKKyFNMllgvrehY2Ji7rmkze+vVha626d/ce3ri36LvXPb1m9AxXZRM2FTbgLla1E5e7cveFd3/4kz/58++889fvMaPB1qePUETKUr74pS9++Stffvfdd9//4L3I2K8bhD9WzqTWWt0rE8HsXEohIjT7IgKQNA5Zh4i2bTdTkQW0DbPy6hU8zgLxGPLo0P6smFmttfeKh0DvXrf99etPHh4etuu193agFf8d4yCKPjM3JCIpE0RHluTkoGROEqI+6pdZWIZWJVPnIDSRGu3G8OCdo1+fTHcSRNSc9ew4iAiAKelQ5abe9JpZhjpJZKogbEwMhdhomhezadg4jusV3SATgy+TKTFl5bxen6CIET3zlHEFW2sRefi9wJCE3oQTUxUiJSKoTsgUQNkkqD9ThkDjS1TEw/4GFWwI0FAllIiSmU/riWiIL1AuMG3W9fT4+Nh7X9eFiDKyZ58agSN7gW5ny7IQEY1EAKtqbZWSDg0xMgpY2/vOLKfzudUdsw6ylJmFR4TDPsbTtMizFnu6YgHpZjNDL0GGpZQIbkpmGM2pthoSw3TOIkaRGe77vp9OJ0g8UG0OljTU7dPplBNjXUqBdszoWsYiwqfTqXf3AVGgMbFkKoNojid4PU+hfEi3Y04qRJ9mZkl83XZAGQalIbJHm00GKTJI2COIXUTHmMAGmNl6B0RlijIiKossOfy5w0nNIvbMB885SZToec4zMzErZDlFMzcuU7eakArY3hlcFExgGSBmiLnNrMAxClfmaT3FqMmwWccw5OnBZI/BHoE01nvH75rTfvS9nFdKkwlCdmYQ87KuRNR6QyE/MzvKO0aSZRAYaBK9mXlZwQHvwz8Lr2VmSALFkJHUn/epIECauXccCT09PRLxMFNPgjk+CqwVEYXY1VqPjFYbC5vqYtZ7h2XezJZl2a7b0aGRKPswPnMpaLvXPVyYy7JEpHfHgFvRyUhxaJfraa17rbUm0VLKspTWcMZRiunoXBo4pMzsvUGgj8mAbq2BZnScC4Zlw/wEHoT4xW7pjBagEQeU2j1a6zIDq6y2mpN97+51rxhZOH/nfWekf5i599ESk4Uj02N+pupeNwBkzExVMlMZZQcszCS8bTVz51loYqoswkS1dSjq/txY1d3r9bq599766XTCfnW9br13EYZx+eH1g6iq6txOZZI1jkUj27Y9PDzg+B8fH1FwcH16oomrzsyIVLny9CxH5Dz35waVL/gZTETJRNdrZuI2jX6JOYHhlHlwIXJuRUSUOZoZeMRB5OA3sT85uucJrM5TyZUItJH0nByQ2a5QUpTEKDql0xuHyd3jk09ev/05ffvtt4koiYvZ/f39+XwJD+JkTuIzJzMxUgL7tpmZmmZS7717x01KVY8dCTMQqVaeFnX5BQEaBnBTRYJQREpGhkdv+3bdmxPJRKM8l0I0p4+f6J33Xn/v3/713/3Kq1evLku/LmqLqQmpJiBkPbiHMGsSu7uaMYPFBKLXYN30PtBVA7fk7pHgpMy+CkFBwhxiS7mQ96yt1fzzb716++mmQtziFre4xWcublv/LW5xi1t8JuIv/uIP4yk99P7u7tX95al/lO1sa1HIM5nMolIyQ5isiAYZEZtSEnn3vXlv+/W6b9da99679x7eGVpqOFGKAAytamqLWimlLCbFykXWVz9/3X/87kff+e47P/vZxyI0GRZvxLIsX/3qV7/85d+8u9x997vf++m77277tm8bEXCDEhn7Xt07RQ41M8cTJgy7RAR5qPtws7bWUIgNSq+olrISZfc9vNN0ovHw+UbvvtcNhk0i8t6vT9fHh4fr9nhgZ4nolwAYQoF+LtyeVEjKIJbkRK1vMocw2A7EzBx8aBaHkjw6IQrr+CFHRFKKHHLuUIiTEholBBH3zszAFWSm9+PROkUkk2qrnKQiZTpAW+9EdFpX4H3dXUUOea73DplyfMr0bU0BOpAJgNAWkRFDgIahGM/bB0f4eA6X2YcNnwb1x6deExkELXISBywUn4nCc/xqBT05snsXFuAvwJ5ArySo1SLioxngGGOas4KmGflodoeDVAPYgYCbYGYABDD3MlOHNa9NGYuGf3AUR+dotwhLIxPgrR6gTwgcpvjtqE+HkRyS1nS3zRnJTJS1VlVNBfTDw4MJWQHHMddacWwylv7QiKFj4vOhoEFEw/XCle1AjaRmpg8RNvbKs0Eii6hzr/vgVLs7zTMlIhYO7+MIiT2HmRFnnRG9N2JWFZ+rOBO2/YDocsi4wg4h7+VUYSbIxGhJCrkL9e7Dspf0TGTuLSLVdPaLGwUN0SokS0wh+G2JxiWOxHhOwZQIvFf3HpGYM+7ORO6GIT1kZTjrzYCMyMP73DsoK2NWw5l+6FCYnGjx5oPHkkiroP4AZ0pEdd+FByj8uKb4Rbg6IHiPlAYLJnyOJZ8Zx1ZESFlRUhPBhAUBF55WoJ+xpQAYraatdUBjhho4mNsBq3QxhQCdmaZmZrW2zBARsH1a6xFOxMtSMrL1kZSyYpSQd5squhRwZoZ3ShaV7h3Qc7x3aeu+7632PljbevS+Y96wWjz8kEFxvY5etVhIMlIOPl6TyXNLzRjMaGGOsRFB1c3e+2D5irh36IlYmCqaGd3d1JgZCikPXvcsApr9HZl5tDoIj0hVLcVabWii2NvIraqoqbqP+TC4QwnWAnJDKsJwp+61YdNY1xPgEsKM3ThJSonMrLV17yKChoH42Jd73cRQPNfxYGMBu99Hkz2qtY073dzp8Mfp6pVIgHRyWRZmGhMex/2MgRiOZiKqdU9KOhr3MZs78hBzgEf9gYtAlpUJkuKpQWNF4cRo7ErDOA8DNVZNnxN7HAFSW2bZInn2fjhulhHb9bqu693lIsxBtNcaU/LNzAyX0VsZrKHwCJozAxJtxiCuIIdHM2k3kujMYxZFjA4A4/BpppnGKzET8JJ8XsovvqhkJpMHPXX6yQev//UPfvybd998285ZPY3So1GYpRqLCXFRMWIhFlVTM2KmPu3zMrLbSFzx/ErQescXlmP507GxiIQuS6z0+PTQ6Rsfnh9Lo1vc4ha3uMVnLG4C9C1ucYtbfCYitkUuezzelbKsxpuW0HUjPZfzcrkvRYWS3L1u2ZtkZHr2Vq+P3lv0nn1v+7Y9PeHJdDw/sZCYLaf11ZlIWFWtsIqZntZS1kWXhbsTKen5hz/6P//sz7/3zo8/vl6bKTdwL/jQoZmI7u/vfv/3/97Xv/51d//www/ff/8DWMxYxB+fMtM9fHS/oePJysySaK8NOg7clIeFsPfOTOGx10rMVsrpdEbzq94qC5/XE1GGO6QrYQny1uq2bSISHk9PT73uPjpZvXigy1+iic5UGmZ1LI8fDlmZBk83OSk9A497RCTEnIz/iGg8fwcnZLb5ER7d3zR/wbAMP2BEUMIyKeI6PX142Xj29t6ZKEXCYbalVivkK5BnoYVBEYAwejAiDpGLiCChQh6cDIrhosIhXa9XGBKfmxbWCsns/v7+QHmMYYNgNJ6ySVE33bsAtts70hLLslASGtzRRFJk5l53MzufTjFUeBdWCLvQMlQVYuX5fIE1G0dCRKWUwd51R2IjMtD+S1UjEqIMGNm1Vli813Wtda+1ns9nEdn3Hf7T7t2nvFusiMq2bdq1lBIZrfW6befzGX58KNrruvbu2/YAJEVrlVhE8dujtrrUwiww0oYGRrK1dj4tKsLM1+sWMdyyR2IgIpdlcB4OuTMigH2AS7SUhSj3fccqL2Xpve+1wmj/9PTovTHz6XR299pq31spepo4l947cC6lLDS0b2U5iM8yMb4BIAacyAFcr5iwEHpXRrIKJVHGwaWNDMrRwispuzdmLmUkAHJI5xwZOYyEEKAhF/Kyrr231tqBIXbkZ7wXs8MMSzBjMiVlb52SrMBNPPINxczda637vq/rOqEuB7x7OG0jIonwyVh3GGERNdPr9To0wTe9wDJ5O9g0h/aXsW27FTufTkzUe79er+uyDIlzHlhEtNZB0X14fIR7sTekiwQZAsiCRJTukGoTsGBmiMJDlJzIXWEuS8FFad6ZuZi1MVsG0QXb6bIUZKXcAxwNd9/2RkmmmkS976DcIFvDLPvDE8YNSIC9deySmdl6y207sg3FzCM/ef2AnV9V9tpr89Zaa71131szVR7QewIxXIX32iKzqMbs9obegd59VIqIZGZtTSZcBfk9D8dki6xMpKa1NuQ4gYl2D6jVWGhQO5kZkKjaWjFjFo9crIiOFILOVJBPsnNR7d1b7yYv+ssyx+g5GhGBBpcdTnAcMxEU5Nm9MzKzlCUy9roTsYq0FjDerstKTEF83bbrzshJMFProPdnKSWIvDUiIeLaHACgGNbhoJHZikgxVeahS7ZaI0aKmUXMdHZoSBVQmIdNXyOZqfUQHg11PcLrwOyY2fyKANLw810znURItWBb0DnrKCg8vXlKPuvO854L2TwikUwiovCwYqRc646jrb1Hhg79OmHTLqW06Ek8wGH5rK57b0+PD0lZyurJW62t9UgqpRBFRmS6ipgV9+juvXWe+YHjtsgs2HXHjqHKTLWOWw/2yZj5jF8MUUEmjCkZbWI7phJOXQ5oGGcSUSP66Yev/7ztf+ftS6n3F99WY6OMtquGFVlPq9jKvIAODgoPMfcecGsftDA64GAHLYRF34zM7L3aspgt1xqn0/rOz37+sLdzyH/7j/7hf/5f/4//H74w3eIWt7jFLX5N4iZA3+IWt7jFr398+9v/JCLzo1dvff5yXrg+fSLZz6udlkVUetvDOby361a3x6i7plN4RO9wV3GKt2iNooM9LMqiRWwty2k5X8rljtRYlUWZkigko7e+bdv2+JRUlvPn/uW3/+yP//mfvH669qAQOigUh6eKiE+n8+/+7jdPp/Xdd3/68PBQ6+h+xhR4qQgnKToaoTjX8QDJTIxHYzJTPBjjoQiMjojQpcDshN5fpVgpysxAheL5ClY14liX5XK5a61dn54OmelX0bV91gsfDGgelGEaZOfR8otnf6nhlx5kaJrPfcPwhf8dEOg3MBvD8iUYDchwNJmY6LhERPCdmenzvx1V1kREFO7ErKqn0xmWK3zuuiwHDBQyBw78YBbTlHJ4Ahlgl2NGwbse1JRh6NPhzhaRUsoUqYeCc4wg1IhEnzQfw5VEwrwsS0b01jLQrjC6OyVBjYWjkDKvmfCL7a2aGIi9hykVz9dADWQmys/XdSVKdKWCOgPNure+5cb41TRAATy4Cj0zr9crVPe9VhmE44CoAZ0dfAZigrI/SMStATL79PQEJ76IPD09zYQK+j1J79E9RMVU1fT1vkfAAolRQVspqvuGyXTUSKOKf+YDIuIE4ypqqQ+THYx1qgoXdkSwSkTU2mAo9t5zThJ4codjmsKD0fkNqgoK8LdtUxEVCeLwiAprKotojA6SbmZWyrZt0O9MTXiwEbAF4GKpByQPiCB9HMlQhnrrY26OH9JzbofaMPFSElEFXQIdIKHiDcRM8OTAwMcnqpkx1GESSjqYHuG++7NsR6Nh4yA84OdmNgTl4eB/ntg+zkVfLtsjQzBexoTJOXy4o8edoNEcjvB0PsuEHmBZjTyNYrlR9ZZwztrA4DwzzrHERNy9hwuPVo6+OzHZYu7OTlaGdIbzEhFNZWErRSF2Y86ILuuSmeHo88ksAQHRVIMF+um4LEnEpKpMnJlJKTpaHCYle/LoYUiZPSJ42pSHQ32c4LOkJyJmZYGyD0CFKAsDTk1EJYmIlmWJgRIao0oLEdFRE4A6Bnrhu1cCCUfwE/e+rMu6rmbo0hm4fNjcYrjFnxOX67oyC9pdArgjInANwxeMFScii5qbLxEw7Oe01eOMVA9PN3NWYlpKSaLIFFXo0VYKNHcAjtb1BGJvEqkqq0yUNupFInNAoI5TxhlEd7XhEw8J9tHfksYLSVharZ24lMKj6sDnLj0UT9xDMbiwz2MYcWONCBKhCJjoc6r2rXXQcmqruFUd4ymzTQOulHDPkdkaV8oHK4iGkDx3eJ6JVppmdg9Xc49hv/aMYxAI5HRmUWMxQkfTMWWPXYVb63y9Xi73Svx4fcJ9LaIzEVEwcyQBCzOyWRga94wIFpzWGKIkUfGIASuhPG59DGrZ4YCe2/zzX5GlTmbmspiUU2vdvWeOked5Aw2iq+fPn/o77/38LYuvvFqScpVUVRKOpOu2i7gYvgHiOxIFhm1ay48tFAMeY1NLwS2Vn/3nxCRMZVmsLK3lLqvXlswq5Rvf/Un+EtVkt7jFLW5xi791cROgb3GLW9ziMxA79ZUXzbvTulDbH36WvheOQuRt26szc29937a2b16rRKfB8QPpQpVSVIueVYuIJotYsbIuZSnrSU8nEk0RIs7o0bu3re7btl0fH68tNHX/s7/4N3/+f3z3urcgjnyjfx+qkC+Xy5e++MWvfOUrj09PH3z4QWYsyzqNX5STGGCUsH3iKdHdxZRZzEp4wsQaGeEdrrZRT83UJyo3IsIDogyzZAQlZcbgJosSJzOJ6sPr19cDkvArCMYjLsR0piEnEwnLoUcTw97MoykhDcMVj+LkqcUOuZmOauiDzjFqjnkIWUKU0ICJKCNEVYRFKGNQMoiIeEi9qCUnSlUVYsqsSczwbGpmHk6xo4fb0dWKiCCtHnoxHwcBCxWx6tDeRSRzyOiosya4XCebWNWOqm38a07YQlISRybK2EUgnouYWW+tt6F9MwyrAwaSMHUOuzcxjK5BIhw8n5Yzg5KYZN/2yCxmcAGXYr1nZnr36aqWJG4OJi9gptl7691luPygvcL5l9lAckj8Kz/DkXMajZl6r0RAPFMSpGcEPohp9OkionVdM6K1Ks5UiqmGx8ECzggFalS4tUaUpoaOfJEEHTMm3SWHlurzd/nk0h5SiR9Dmkm9NZ4ZhUPWwXrMIX4Nhy+yHNgtmLnWyiyqRsLpER7CnCQJbi10MCIiaq2DBIIfu3cRHXN4HGTC8S+jFICmcMZBGR486wmGRDWMzxMIkjl9hQMgjtRLRFAkEZsY5g/kWfwizCMVEVYmNhWabFbPYWQuxbzj3KSUomqtVT6Q5Ul99kVUkcNMijfmQKjDMX0AN8jMIpN7U1UB+TcyKddlgcTTW1eT0+nUWw/3TMLGGRMnDQ84+6Chq4iH9+6ophdVysDGUVvrvevsMTjb063de0YIzMKHfT7TMiH4soyEDTOpmqiEe621lCIsnkExQEBHnomZCxVcyiP/ZPPZZNDyZWx2SDL5GPMh3RKRio1tk0hFQBnKMjZNJopxaSRG99PAfQH5gMx4IfqPqYUldoizUHVjcPMhMRsl1cwiYmai0FLb8IaKCI9ueB7hA2KDTo+cSZGOO0Ephm08OcNDCPZ/KWbo8ob0WGSMSghVJCrG3Y0I+KxlWXpGZNjwJtNSighY586cp3VFuQNmLFrIEpGoOpYAUDO41Q4XPIXHEO+FWQZMI0e2VLHYRa3uNSJkGm3nIDD6+oLeg1vTvBHovCFm5oAvsUiSE0dwTH8xT+CFEJYiC08wBhEfsisRE9KZODdUPGTO2yOWy9gjhFlZiCgEO6AkESoAmHn6fQV0rJj7nphjZDkyKSYPGqvMW2uZIaqmYxRKMSLQKTiTwMdXFnRcRD9JmjnawdnA6NlYCIoCkdHKb+5dz19Fcuazh6A/VkRmcpqaikZuAPE8v4MISZgW9FjzR+998vbJPvfWvXEWy1NZFmWRREWLjh6/iZsFJ7EO1ldOxAaSTN2HuD6vgObsXRyZxGSmZiZiHuTLffSWWerS/+P/6X//s3/w79O/+B7d4ha3uMUtPhtxE6BvcYtb3OLXPL797X9MdafXa56Fw2P/+fbxe9keJaurRI/WQsRSjElXUV5LBkdqZHqkmFpZRKWUsq7rsl50WfFAyBlRa4bH9ujeMp0ye9t73TrKoD3W5fLwyfX7P/rxj/76vY8e9h4cykEc1OfzE2WSJP3ON377W9/61vl8+ejjj/e6/8Zv/OZbn2t7bcLs3bdtExU1naW6XPfq7qJKTCxystU9sqeZjYdHIg9vrS+liGptFSxD915r3WtCGenujMc2ncJHuoe33l9/8snrT15H7xREJP831OpPx99k5ZmEDdSSBzNzMo3WQIzCXh56HydRhhAJCUsmZdB0/SUFnFrDCofDxe+AdRcagypPv9h0jk3qpSosiTSsqTwMtXCZLcsKzZSI8dQLRRWvhMAEO3OrFb/cvSeRsJipTGYxvLo4qlKKu6MDGDOv6xrh+77P7MIUf6bQbGagFtRaI0YfKsigy7Ks6zqK0BkpA46AQZ7IMyOFeV1W9E6MTHfvrVsppoqaejULd81crCxLEdEGRVVk6K6Rqmwkp9O6FBt190x4NCciFTmdz8J8vV6jFGbCuZ/XtfWGc4RqmagjiFjWNTNabaUMQsKr+1cQ6+F98xiMFOhBsAdCmEagd9/d3R3gGMuywKoL4S8j7u/eFoHNvGXm6XQCFOJ8PvFwFLbDYA5fs4jAut5au16vp9OplBKRkKrhAH1GQBBkvnQzFTEzFslId+ejgaRHUi6lADOCtooUVEph4da7zKSIe3gPnvCBOUNJhi9UklJVUVzf0fFP9LhAQwqcukxoHKZ9aNaQvXI02Ixjmoko5WghyIMY0HrvaiosTGMKmdnB2rbBBwc2iEb5RQ5jLJDWZuaZEJoz0sN7a2VZlmUJH2AHcB6E5QBtD6lLeKrqiKNLG0+f8rA8Jz2rUMK8rGtMLLiqnNYTLjEu3CFLASaTmUdvTCQzmBm03GVdWq2RaarHVPTuvff7z92xcO++BDpSLjnJIVNoW5il9wlPv+OkzPDuTpZ35wuurwPGTVx7hZPduxNTsTK8qN54qlcRYBOnjK6nMZRiLjx2y5GSgQ18XPQIEVXT6E5MopqREZ5B6RGRwpLESTL5IT0H2zqQTsMe9dJFC80UE1SYe+/EXMx6rUN+ZeFEujaIU80ys+7bejotZUA2qndodrXWogbJcNaZDKG/tZbuwilCWDQslCmZwcIqXIpizHVKz1Asl2UlooxASjOZRIuMXVHM7HI6I6vn7sHBzMuymCqmxPDVUialmgozLiWyIxmovxFVUdPIUSuAHEbvzsIwkmMPUwFGY7TyE1FixuqjkX4TVYHH3Dss7DlvXorsGrb9QYZBdcjsFmhq+MDeB1tJZhfIyMjI2dXQ46Ag8yw8yVHdwS8s7THzUTSN7YdD+tiSwNVh4qrSqpIHR48ON3JywsAcH/385+vpdH85bdvOwp/7/Od6923fMwIfDb6QmcW0C8/NkCMzHHhrEpHe+gTEH05iYZbuI/05eCwDZ03dOxEXM6TT2IR5qP9z5ImGbXt8FwiiLeL7P328v7z6u7/3KhfXle4u5a3L6bIWSkciW9E9AYQpEmYxUzWDgO7hrTakpmK6uz0iPAAxr/vWHOMb4dF7hHdqW2G7ZkjGf/eP/uFvff+nf8O3plvc4ha3uMWvYdwE6Fvc4hYe2h31AAAgAElEQVS3+DUP3u9y/VD7V1fW+vi6bR/1/SnaI/tOKpwkQUoLC5OVcjqrWfROIqmaRGwmpXCmsphZJvcGgmNPb9k7eYteve8ZrpLh3nutbfeklCLL8sFH7//P/8sf/+ivf7p7BGmOVj5ob8NMJMQq9tu//Y1vfvN3Hl6/fv36dURqMSNq3YWFjCGCAx0wpSVSCCWAHiyLRYYFJbEwirIzc1mGx+1yd0GvvszFrJiViQam0ZUPSiG8oK3v27Y9Xeu+w1r1y9aJ8vAw0zA+Q42By1loUjjG0+/xN2hmyuMdMvsREckLi/TRI0sEfeoJXaGIacia8tyaDH49ngI0eCZmVlsFwOTwtFLCYzYECCLKzHVdeTzWDilsOHPNRgV9RinFzNBaEHpHJu37DoG1FIuYCiAoCpPRASFWhwVNJn+ZpzMxpoFuHDwdDrJxMNCc80BS0jxrVRPh6/WK4zms33jlgC7kYc/002mFKXVqguP1l8sFZw0tT+exHtfZPZiHp5snTDZmm6alFBCcI1zVULl/fD7+UC4XKIM0LO64wsMud5AciAZ7oZSSGa218/mMMUR7t8vlEhG11mMiQZ2coj8DVQzP+7L0ZVkOSXTM2VlkgL+Of+Khd2OcofAiE0BTuMHSixwt6QJ19UmnU4GHt/WmmrSMiXRc9EP3WZeVJih8rqCpNUfm9M/SaESW0/9PxxzI4QYksHN4Imggf2eMnp6UqWJjak21ZvAfMmH3nAR2iFWhasTkfbDR1wmZWc1wLikpIkspOOajL19EoMQe2ZEc3mHtU787ZvKxIkb/QGZsVocmjomHU4QshPe+rD/AT15ezeMPx26AjWHfNjpOOZNhJV7EbExRSpJSgPeBPp4pcwMRESWbswrb05wPc42TzW6xE/zNvA6FbRqcT7huLAIauNrsHorrSaMIJjzdw8OPpYRue713ETXIcDl61k2kzMhgqaiVMjeWQsIJELBZKWXfd/RFPEZrzOfZr+/u7u7YfwANx0knUWR4OpqOqupSFiRdhGUpZYALkkeq4chlzn0erRdjJAh1bPVJzBwZ7rEsy+FQftE4YdTIABFDzO6O+ZiTGQXG1DgfngUy6J0wg5lEJTMo0lYLd49QFlKCOm9mVrS7906UOfauoctTohBh3IM4CTtqsjILz/wL4agmnUlKKeCGUxK8wc+3PNShiKCV35y6jFIhSrEimSwMO3IQPMJCMe8DhwN6GMwzRURNUZHSvYPZTRERx7ogZrTfzJlfwRxmVSEqSRmZEXvEKGfBteRkiqz7bqal3KFuQpiEyVQEfXqJQoKZrTwP+8wic0SCE0U87uyQ6Z+Tyonx1XiTW4XPwao/Zj5qlaK7MO+c117nbHmefEHUkl5Xf/f19YfvffS1tzQv7PUpwikvTC6UIiSD9iSZkRTMksKMuhnsqqWYGc0iLYjpmalm4bHvO1JVIpzJGeThLbTy8uHj9fVWm/Bf/t7X/vG3fuu/+K/+Cd3iFre4xS0+A3EToG9xi1vc4tc5/vAP//B6jbv6m7aYZlxff0T7a8sBFgYOUkzNFikr2+l0f29lCXc2k7KQSqqSSuxbth6Z9elar5UyM3qmG1NG721vfeeMUpSFk9iTyYqe7kNPP/ngo3/6x//iJx90n+Wfx4MhHIellLvL/Te+8Vtf/cqXv/+DH/zsZz9DrbB7h2kLlZ2oumXmSBi+RFVYJgl0dtJqrXEyC6mYiWih69OTh9+d7pk4IkW4FGbWjGBiFXHvLROKXu8d/tyHh8e67eH9V4DfgHJAzCw4kfGwDQ1ZDrTzQHAQj9JjKE2qxrOEeaoHeLSfJmgIT8JEpO5EWZZFZhX/IWYRUbjDaDYE6Aw4l60MvycdUp4AtJxT5RnP86isP8THodvC5tw7GBqn0+l0Ou37DjwF2ALodPdSDpvi7PBpzg/EidNxqqhel4n6BTcZxw9z7jqqy8fnQLk+FNsjcpIilmU5nt7nkWittbUK7ges1hixeUjjTE+nExGhOWFmllKWZYFb1l80iTrKotESE29xj1IMHJUpMo4Dw5G7+77X8/liZtu2menRmeqwtbbWoBQf7RDXdcXlOHrfQZZdloUm6JZfWHoPs9rRHA9i3Pl8hkINf7SMDnXwyQ4iwbiCzK1WOH+JSDVUDdPvsCTTMeuSInzb9wgvVsyMibsHS6qajKHwqXXyRFKA8cqHdRfi77MArQolJAJt38ZVjpmI8JhtMCcD5phszEz6TBcxmwT1ZCaygff1qYiN9l+grLg7KfC46EzIYB9jzmRm9w5pclkXeJOLGYtQZuudMjvYr3PGRNjeKmYUriys7qUUXO5a62AUDA87loMS0bZdDz06M+soSoDGx8wM0netLcKPdYcrDhEWFQ/btq3rekz+TMJqNXtujIahOBok5mzj2aiJBjivgDbMVBkdCB0GwYEIbB9cl3VdmQ4QhCzL0lpH/QSQLWUpzNR7w4Efl6NVF3FNPZ1OIrrveylmZr11JCnDQaPxzERzgMxw933fSymXy+Xh4QGjzaLE5O5WylJKKYZcEWhMNPktptpq3ff9/v7e1Fpvw8P6Ii2ZPDIeGFWenl9bTRXAZ2ai3l40zaMM7BqZpRQ+kCnwVWdmpCiDIL9YwSZ/5CSImJKP3FcpCwv31uf+zT289U5TSrfZ+rL15t3LUjLJe/cIYSpLabVGuqqEu7fOZgwMN+5aRAQ9P0IkkjSn6zVysOfDHSD50TgBfl53pj5pFTFTdGVdFZUxWEcySzSwPwkzCR2X8jlvQhSUpoWYPANvUZWj4ufojjhyV8yAaZgidde9e+udShFou3Eo+pzJOXsX09zEiEKVmTXTIv4v9t7lSbIkS/M6D9V7zdw9IiuzsruraqS6u3oYGKYRgWGEPQhs2PBPsECEEVjCli0sQWZEWLBh2QsWgAybEWFEEJqZnn7SDfSzqrLrlVlVGRnh4W52r6qec1h8qmoW2QNCd7GAEDubcPcwu3Yfqnrtfuc7v2P7vpHbdTo6KDjIW3NrTL6uCzN7q9Ys3FNeiNnM8crLLbznDqZ0O74p9KSRGvj+PV8SPV89Wh8j6Ys5iMVBVV0kiHJK1poR7rx2PhNd+M/9vUHUiHaiz5/Pf/jJD/kbH0jLb+257qXulb0liaTEQap6WFfcOUgk52XJq6hQULhLSqw9+4AEVRLg41N4MGuvY1iWpEkkEZM5FZeXW/v+j3/yxXN5Vv4bf/SD66l0i1vc4ha3eI/jJkDf4ha3uMX7HB8+rD98tf/1j0WVbXuMcs6ajg8fC3+FyUQodRQyi2TVg6aFB0XTqksz81Mp+/npse1bRHht0ZxZkkK4zI5q6+CQHOlAKXPKL5Yl3b+I5f7P/uz73/7h6fs/sdOOsnmaDq5wAmv2xUcvf/VX/+bXv/7z7u2TP//k81evzUNTAkawok2akbsHhQo3a7XW7nQWqa2Fe0qJupvSUtJ1WVJO4XHeznh+S1+8EU5Mam54RuUgYdYkQw5qoBlu23k7n8+nU63loob+lWVo7i4/4iEjT7tyl6GHFRr1vzA/y8XGOHvQU7eaMRPjaU+Ha4yom+lUhZi1v55giORpTIThN7rpC0/mpda97LCnGSp/RVSFPIASJiIUCDOTqEJoTilNdIa3tm/7sM/yvu/7vo9q6Hh+foZqBukEEue6rufz2XvRdBezrg3OkB25e/qgCTp0tGVZiNg7xLa7dAesOee8bNs5IlLKsOJObAiEM/igZZ7/rsDSpE7DOIyy4ZSyiIBsC1t3DAQB3Gf4UBru7+vLzswgtxKq0SnMLGeJ8H3foSpOWRxqr6ru+1YKWv81SIrY233faejU0CVzXtZ1QSPBeZhzx56enq63PAy+NPtDzj9CjpxnCdtvDWY6Qf5gHE4XQAOcmt7oK2ppSEKUUlptHRGf0nN5dnfi3iNuO+/MhYfTtpQqA5djzQqzphTuzYwoQCcATzk60FcgfLg7w4DckRzh4VAwPHyqOmOI9yPFy2DglcF1AdxDWKAGmhmKLIQFJJOJ1IAVNOe8171ZoyAgNbo/N+Lt8xOsi6VU875ZYnafSqhA8uuKLLM9P7u75oQhh1FXSjkcVvSxxEibE2HkLWSYkbsECPnyemQikaMKEzGbNWYGDAfjIXorTougUip4LCPhEedz95IjdbEsy/l8BsFmzhozN2uqUE4Df51+VY/uPp5FBshf0EgjLcsqaAzIqLHoSHHhzrqPrvFi/OOv1DVuZk26bRsTu/voyimaNGnatq22FnEpmMAQIebWrJSybRsmaTM3GJm3HVwIjI0YNynIwYAbtGpvH5/mjnUADqo6lkxEbVDdsSy4OxYo1S4ouxt5MHHShAXDzNB0D7SZwZKOfiHMzZpHMPNZepPGwebu1zppAjZC9nMQmUGpZGZqZtUaOh+6m1RlIhupxGotPJoZhNDzfk6qTHx6eiIiYa6Gjqxaat1rZQoWIeJWWzVL6BfoZqUs68qqWDFAavCgZs7VVGkOFRoJwoiotbX2HEDpqBCLObVqzJxSBgK+NtMkzBJhcONyb+FgJKqiTpSThDONVpxJUzCbdVT4XOgiKLxt55pEkuqSD82aWxVW0gGp6HniIIokHNThJMosKi3MhZJKFXYhjr7MdHY2YB37/uaLLz786KPD4dianc7b6by1ZkHcxsTsyYHew7Gn6nCvGXeNfge01lLKy5prbUw4LdVav02IykiwMYHjH+4RwnxY11LKvu3rspi7aA585+nfZlh7D+IwosdT+eQHr375qx9ouotWtt0en87RSlY+JA03YTnnilyaE6WUc156CspMl0VVmUhUQPvuXWU1EbGZpaw557QY3OsiIpol5eO6/sJHH2z7T6nZv/Hf//bv/Wvfon/6nb/qd6xb3OIWt7jF/2/iJkDf4ha3uMX7HGviX/nayzXb/bKwEemS03p3fycSQeZhzEHCzY2cpZl4ZWoN2pI3cnOr1vbt+anVnSnIgpxERHImJeEkObFqFqa06PGONbNmXVZe7p8r//4ffu/3//CTx3Pv3wQuI3d9KNCZ58MPv/K3//a/8vBw/+bxzePj2+fnkxOlpCxKJLU1M2cWQ/Ws8EDmhggH/HTM3t24DkmitmbutdXT6YSq/20vQsYMyY9UxZoRuThqyS3waNva6XQ6n0617DEgkhck5F82+GLreadZoIxqYu4V/9dmXRqqMkqXoxe4xnilzMJr7438LqQGUE08AkjpXmvfVZ5O9pyGKLzForuoiDqyA2xpAvLTfdi3CUwPeE5bM+auT0WAGszXVlNVxVXGxZrCzQDydnMrgAkQPVHrzQN924WSWml8fAx6Jg2Reupu0SvtqTUbrkkyY0h72EkepfTTzBuXvkkdL9Bag1MSqllExT5AR4PM3ZoBTYBfzWyCqodWbjwskENMByijuxenBRWsTxk0kqHCKxGVUmqtkNFxuoh4KM5QqcysgzVwQmiASmgIzRCsry3PrRmGG/zj01iNs0SDmwyvqwhDOcK5NXMKyjlHb27Wkx+11IhY1tVaa60FkeyiKrVUjxDVnBIzl+5vZWQ75q5iuHF38vZ2iywsogPfgVlOgkEV0TNC0V2EQwvnGCXqAxKN/oqgJVBMDobIFAppzEq4LStSPqpWq0doa30qmCXVoNj3Yt6YGbCDZg0ZJMiXqtrXz9E31dxpJCHCvdaaehUCt1qb2RqHGM5lyJT7XvAz1rpa20Ra01UBPsTiUYgf+164Z6HUzFozAMe/NCow2fGWq+10dAxc8swc4WYu0rkf2763MQu4a83ozDccyhMzMlYtrKuYSmaeVE3EsNj2WcxoYTrbpfYueQx0AwR39Nu7wq0Qq4gmNeRIwPQgHowm3c5ba4241x/ANs6EwUNwQ2MpqM0NquU4hyCuDH8zBOjRs87dBuAI+xboaKequ3pEc5vjGafUzIDvxQlv1qSrw13oDECoibSzz/tRi3RQcreud12yC9C4N+B+px3uEVAhca8ERwIiYwVD/IpqjImBpdcjukE6PGkiorIXgp7Y97OXvwxMP7fWKKaU7LW1ai4qzQyMYVBwPLyN+psBDScREYV12s1cJSG/2qoRU61NVXLOZS/NLMJTUmIqpYhqBxZht82ZcbDcx6q7e2CGmrXrtCsNw364m6akyiKtAYjfwex9Gemwl9Ha1KOPT+Faa6sNIvu4rTNdnVaiaK2dT6f7h4f1sOKc19YiNqLJCUemU/oCGAC5KK419eyzDHnXmVstZGa4uJi8uFrsgI9JSho92+NBxNLvnuZeW4sIzclqhDlhBSS0PEbfSd4tXj1uP/ni+Rtfufv6V76a2EtrGkrEIokZSB8RSREc7hFs1jMsrTUBx38suTRI0z2fbbYsKeXEIiRM3RudNGXJB+OF3c3qf/13/81v/slnf+HL0y1ucYtb3OI9jJsAfYtb3OIW7238k3/436SFVdrHH35wp7LePUS4CKsqMVm0fT+bt+pt37dWLBotKVPQtm1u5uGtFeXIKlYbOSkzXMxOjCZWpLqsh7weaFloPdDdHZFEiDU+7fHjH7/5n/7n3/zN3/mDRgFPr4fzQLLi0S0Jf/zxR3/n7/yrn332408//RQ99lptzZpqSimj/j0lQYV8SmlZcvhSW4P6KaJ4ZIM/CBZgPL+5eXgc74/Lum7bHk6wyuWUlpS37YSWcbAQQWcN9lZrrSXcuuD7swcPrXkYnKdkfMUCpfmXSTEQnrZNHy2SQiSIyCK60DwgEnhq7VzozkMgGWIuEYmIq1JX1KOreDhX4UMVR6c2pqFSt9aEZVky3LU7gAApuzX3rix3/HRrUMpg8Zru3ZwXES5ln0qTXdnBoERM325EiGj3UEZAPnYPVaA2YvBbKToVgYA5FpFlWVtr23aG8DRFXqhJ8Jaa2VTAIfnBYTr9yLXW0+l0f3+/LGtKvG0bzKHMXc5urZVS7+6OQ+ZrV9eZc85EtO87zvmyrNCJ4FMuZS8lg5Ht7mj9h3fB8Xo6ne7vH9ZV8PO27Xd3d/Bx11qZBZuC7RrchnnqpnA/j4WIoGAOz+miCiG+N9cCuCOunLOQOzFIUUaP0wuCgYii0n8mDCDin0/nZm0pe0qJiPd9N4ACVERERXciRz9DvspShCPZgZSAiMxMjyYgj32kZhRAnpm+GYzXi+4JAZr6SJbohQQ9Z4Dto2tixOxhSEFk1t3NUKysNfTgw+SEMRxrhFOUng6R4HDqGqGIskpOitQXkhvTayyirL04w81AbWai2ZwwwnlkAph5WZbWWikNrBgzb81yzofDCh/imCOMpnmgxLbWnp6ecs6HwyHnhagCIz7mVFe1YnRKnEUDXadjIiIzJH7ATJcpT2/bJmitOSz2s4CgNSNi5I0wSokIxGp3b8YpJRV1dWb28NYa5nLXBLu3njs33G3wXiRwScU9iF2GquZADTSzUnbv9Qd99iGxVPbSbdEi7vH8fIpBucGH4hP3bUdPt+7pJjazwXK6pPQCOF0RVT2fN2a+uztOMgyPqgJzbwHIu15kSeoZu+Ph0Mc5MwWZowqBUNoSRDbJD0RzV3ko12YNeUdm3kvtnBBmFalecYNQVY+oFdZ7NvekmlM+bZuHq6i7B0Ua4xyclp6Ei+Ag83NQqAjyjsuyhPu+FxZW1ZySjVuJm4d7zomYmxmfz9imihBx2XcRWZZlNs2bNxckTaF9W+vAa+2Gd2pmaBKw78XdRUU4gBLWlFJOTjGQxGFmpZYlLykl804yka41AzA2xhYytYACcaEg80upCmYrxjl8yjKWcTOUqmiv7UCtiXnvcUw9xTg48xTupfh2Puec1/UgIkJcS68tmIsb7pgRFKO58EUuvwqQsogCPGhDM0MkUXo6xEXIQ2qr/W7I7B6n/ayj10IQcMyNfKrmDKIKh6skpzg1//NPf/oLL9d/6V/456g8n9+8WtJ6t+jdojmrMMMoEES1GvYV67+IOHIXMRsrhrnXBnkaZTqZhatVltE/WoSZ83LQu6+ctlpJQvRP//rP/71//1//u3//H9EtbnGLW9zivY6bAH2LW9ziFu9tsEQrVR+W9aDcnrf9DTtaJXXchHlzchfomLKkJFSJIqsZmZkHE7MGJ1kXUU05o9/duqzLcc3rojKaeylF7Pb67bbX0ojyy09++MXv/P6ffvvPvvv4+q3GRdAcNMIgopT0V771S7/8S7/k7q8+f/XjH//EzO7u7l6ktO9bEOTmZWgoGV3v8cCj44k9dYddO+SERlUEWKVZxIE/fAlp6W7NMD+mnIUlwkUWs34fDIfy+Fz23Zqh1TwRFOK46MR/2bj2e88/QXpzIfaO5RiqCHWvWzc48/UzI7Ogb2OvdScGyZuIiKZJEM/DdHEkdQF7bK/vjfaScB/Fx8SAIQQar6FFVVfwVbW1jigtpaKQNgPLizZ3wjKKoOOKKYGfS6nMNPzOBObGNBimlICKTknxmpxzBJnNLnwc4bUazMJ81V3Qrvrjufu+F0jhE4Y7yr2rmaWUxx46EZVS9r10eix8u8NYDXV437dBpBVs8/n5WXvXQd62La6CiGDfLqUMxZ+ZqdaCF0wf95SD4QyF5GRmgHWY2fl82rbz9BefzyfsNtSufd+GjU5x7KjWnwSPnPP5fIbLFYe/bRszHw6HiNj37XzeRBgiNQ4qIkR1ycvpdG6t1Vpz7q0Op7qNjUfEtu3Y4NTp4K7NeSEiWJ5ptGccggpFkDAtOfcLSiHMwt1wPfzonZZA/fIOdZnIvRHP/nU9sxKXrA2pSHQX69wvOExZVTTJsOcFcYzsDIYRaS/vpz5rYK0Ov4B7mYU5pYwLJCrKSh3zHTkvF/U8Iuc8uoMG2pqmwdJ1M1hHxxIYEOAiAuUdYEBPu+i8su5OxKqCi4jLOmfB/Pnh4YUqeprZ8XhQ/QpE8IhY15WItm07Ho/4CH6neyeWCF6WftFp1ByMnb18EE4u5Kecs7VOkMD/QlkeF5FGi0EadtFY8uIREa6iITGENizIklJyzzgyVBV0r3EEM2PKDDgvixymgE7d6t5H4xS7p6Y3HNY9S4TMhAAqMcfZkNd7eoIJ/dz2ZnZBuvNccOiqg6iIZOoyPxOD+S69nyHXUsOjtZZTZubaW4xySt0bSwRb6dBMeTD3Jfq9QJA4dJupu6BKvbECM7fmRCF9ySc0PNhraW79tAy09GC09ERUgJuhEGHDg0RUNVMEk6zLAfcRLClJtdSac1LtNvCkCeeqDxuKlFPPOxGJc1CklITFzChcmBVTSTA/WkoLLiuj9633jnu4panKuqJ4gYZ+qR4eHDktKgm9A5VilEaEMlk4MyVNuPNKrwTqjCQsLZfEUjBROAkxKWYrJFqRlImZLZg1KyuJG1dyAQuGwsitu3678ZfP2y56Smm5v7tLmh8fH4N4Xdc2snxLzprULQZHXjzCWpukHRrZlIhAj0181WFhIhlaL+uSmJmFRNmDgiMlxUKHu1RDWwIh0RRE4UbuEYTTwMTmzhRO9JM35bufPf/g1elBmwR5dG6SCKUkSROm9HpYkDK8vvMFeDv9XuEWgY9Ftt0jam3nbYM9XnoJQrO6b29flyZNF87akme9iRK3uMUtbvH+x22tv8UtbnGL9zP+5B/8g6fYWnYhL9vJ6pu2vRVzsubWvDU3i3AXxhNhSkmVvDW0GBKwX4lJEmvmvGrKKaVwF+F1PeiSSLiUXcKyUCu7lZOd3z6fym4qd/yd73znH//j3/jBDz49n3eiq96DeJwOYqak8ovf/OY3vv71fd/fPD4+Pz/lnFUz2ka5uwgvKRFRM1MRFYGTy9yPh9U9zts5pcRMjRzSrQz3rDVm5rws7uZuSZNZC4/DITFzaxQB7xWEV2KiZ4/z+WzNIOGOMv+f8VLw3AbErPFrDCNV8CAJQPyVkCng0JDTmKQ3cfReYs0RvWcgDNE+xdm4Eq87AmIeiIczcWjX8S+fAFMYHj4hYqAKuP/sNMARFMQi4U6E6uBucCPqjQHhPeRL7XbjYc51D1RSE3UK7bRhivAUgrm7KRtRzGaAeNe1MZOmvDTclyKSco4hm8LIBjGoNZt8BjzPn07nw+GwLA77Niqa4YYE67m1JqIpqUiUUvZ9SymjNyBgGiICGzj8m9iH6CCOyUzouvaU/Mxs27bWGpRu/GXgXnjfCygBUDZb66ZX0FHcZi6h4iJDpuzHPngawC9M/V2GlNlaA5/EzNZ1NTMAi5OqirQGuvQOu3HXcQN16LNLJLAhklQhKg7ltONWINFOkAhhz0EzT9qpzePCQakU0Tl1kZ8JAql55FQcZe+whQ6/7hWGA2IlnPF96kb/gTujoIsmcxL25qUDeNP3amaLYhQqMFF4gNkaQR1awEQc3VKamDrFPIiAk6bLPnYQjndzpehQOTGYk2qzRl3T6Yskxsm0wV4rzjizU/SMAe4QEajM7g7is6pORkE3uo63g/SC1Mv1JKLR6y8GmoZGNisG13jOvghSjX4yPQDW0OvepMzC6uZgcmMuqCiheJ8lLmkkn8jm4W8N7imDmO09VYRVwRdCrYeIoO1hX8I8+jIW7u61tjkGpC9Z49IwOCFBwSMdRuiGh6weVmRYU6fvGxAbnBBRZZEwoyvmfkxaxfiQAQ/qY20kWHrVyLjiSHainaYwc7iP+hvhgZOJMeiZSEWpy8j9FiAo/XH07CWehOKeWSG0vCXuJJOJTOAxBUSEei5UEtqZMolKeAQ59RIcUe2ta2E1HkSRzmni2S6SKKmG8Myl9eMd2GLJybxgD3GeNfA+qPCk0ndQU8/K9AQsMRMrwz0tzByjvgi9QYmZQ1g4aeqpLACOuGcLtF8hZhaKuDDmk87Dwa1bZ5NYFZIItEBuxBHBFB7UGSp9tSEiVJY8PLRlWdd1ySkF8bIsyd3dm7smFRYKnwk6d1cREJD4ygrdR5oIvguh7sGsH9I0bquqdNJL4k7oYqE+V5hDcmbmWj24gwy8/IwAACAASURBVGwwKCLcKZzocWs/en3+zqevvvmV5aM1BVV3czJ3cndS9jAP0EIuaXIhip7EoggGUCQzs2hEqCig86W1w350fMdyB9q8ln03lqxnl6a2LIdq9p//B//2f/hf/A90i1vc4ha3eH/jJkDf4ha3uMX7GduhPmyHx/UpCb15/Rntj2zn5JGZF1U0Ljfvjzeak6YUItWLm6no3fFwON6l9Y5TJkm03hEr1xZWww1EhdP2/PjmTVb+8OXD28dX++lttL06Gx9E6ief/OA3/ulv/fSLxxZh1FuBvdPpPEhZvvb1r331qx+9efN4Pp9Z5KOPXp63/en5eUAG7aiaUlIQHkrl3KkCtK7CzEFmDfoPzEA+oLLTOjf6RUVrNdxzVoXXBrpq9woHB9W9PD89Y4NjX382+ZnnP8NgCeKkDMWn/zMeq6nDAYCupKFhjAe+CSRg8uAg7cCM2TWLu1oh80T3MzB3BXpQ0m6Vm8+7EUN0uzpozh0hDfoBDTwrMTdrMUQZimiDTTmV0NwfeutUviIiohNOp/vSLi3yZIqSKKWHPIrnefiLa63btuFB/cJtuHB+udZ6Op/hcBzHT601ETdr07aJ4eFuEFuZO1i8468HzTnnpZR923zIatB2mwibQQHkUqqZHQ4rxtu27SJ8d3eP7TNfK3oE0ZmImMU95idGeGvGzDnn2WjR3Utpvdw+6b7txHw8HMbUQMfF1NtDueecI+Lp6Uk1pZTgIo9hSj2dThiAx+Ox1lpri9hSSvf396UWN9v3PefleDzCil5rPRwOnQxubXjxUE2OVnUuXWpSNwt3SSmYggKclnVdmcjMSyk5JxVVEQ8Pp9STCoShL/B5Ejye4RyDhNDlPuJBpnGHYzWuDLbcu4ddb8K7vXk4eWksBDRePCAeNDWgjsRFjToMs+YTWFxKEWYVsdZlLvQytdpwffdSiSJpmrxmcEFyTnC4e4SKrCl3Na276cWHAvr4+DYGbBcnupSylyLj17FZn78iqQDv5Gw7SUTPz6eR/pGU9OnpCadnduDE+ceVHdOTkGmYJl9mRjFB6uUOnbMfwzGtqsKdzDuYM7lr4g6fsgxue5d3RZW647vDQMpezA2UcEwBYhqi89SGpzW+37PmAuJQ9ESAYUAzAIpg4YjGLABhx6AARwRKJVQ1oJsPHsPsdQi1N4aMvuSMrKeMc87MSURVQxUGcGhr+77j6izrgguBa73kjB3e9+Ju65IPh4OoPj8/E9GSFoiMHVnA3HtCJlXtvQdn0sKEieKwHoIIiSJ3i/D7+ztVPZ9PGNHdSCvwHYf0KcMibEw+2zCMDpatmagoca0F6U0WpIPM3FjkcDhYa2625sUjrBmDEDwiqQ5+Mdp52rKuRDpSVpxSYtKIqK2KCFJ5mIY60oqYwUoYgRzeSRoSfbnAOJgfOgtB+lLgaLXXGdbEPAsyuEOZKzHnlL3nU9wGgQoI8euvKUFBNhJXSH8RhQupkDs5vNdM3rtERARZmEerrbXmTnDBY6Yvy0JEzb222mozcxHF7eB6dk8QP25wy7q0CihNGpigQKIL+cu+uqqmlCLYPZCkd/flsBIFUsu1cm2F3v0yAOnYiCrR69P5j77zvYe/8Y2vfeXD2N5Uq1uxRC7Mm4qZoQxgfM0YF6uXudCMZT0s68HMG4uHqeq65MPxoJpEtLUqzFk1yJvH1vjxXD57PG3mbykdlW5xi1vc4hbvd9wE6Fvc4ha3eA8j4j/59u89fnE6HlSP2erT1spGVtOySs4hAgogc5Aqp5yWrCkxS75rFJFU87KkJXMwOYU3Ludwt7KT1bBaa93LVvZdagnmZ9vKfmq1EvHx7mWlwyefff7J9z770Y8ft92DNIaZjMJ7/3imu+Ph537uo4+/+pFq+tGPPnv16vXbx6dtK6XWfS8enXJo7inn8Ki1uduSMjSXbSuiSkx72dwN8FliSklTyiml817C/XgUUWUSs2LGQVJbNLPWGkCTqimJuvnj28fn03OzGrNO92c2Pw9PGNNQleAOHgI0RB5RFjzIEU8BegjWfQNQqLs9S0Q4SAiI3S7aTqFmynF4Yofy1j1qaF1FocJ4Yp7vnbY10AAI/bVEHK3ZWn+K7lY3uJvdoXtCv8Nj6PF4jMGZJaJlWaL3l5OhW9HFHjuMotj7ZcnzvEApLqVAlJnlye6xLJmG21pEDoeDd5B011y6iv5uS0BIPFfqW1x5qDuxV4RHysJVdV0PMCCPhorzopI7WllqFxMHXvbFi5fzkhGRu00x3XtvtyCi+/v7oZB2o72qQhCU7h/uzd/mTi55wSnC/tfaQK6eGGhIGOu6qqqIttag3UDL3vcd2A0RKaXmXEUUqI2jH3D4OS+qUuuCjwbzF+cDpwVi7oBdwLDPcBPSMGZT912yiMJLfO8+tFY4QGmI8oSRidOL+RHdcX851TzyMSjPJwzkefYu7Qb7jIkIbzYMoO8OshhFDVdYHb5YeiMiyIfp2L3rpMTE5Gj5Jdq8mZlbEAUPWyIF5VwpqLdKc6+1pUUV9RmtCVZd4aTJr1rYEXPHb4cvS+6HOUJVD4eDivJoeIacDfQm6t7DOqcbOlL2ZUUYo5R7O80+9Yhotr4ciGEfOHUDJHmuPXNZwXuheY3OgUzUobTuLsZEBOF1eqWHAP1OGYiM9BvQEOu6UNCyZFyT7posJQ/R9sIkGQgmZhYdsxgdVqkvksyMJQvsAlUFxMnM3ByaOBrQDcGZKXjObgd3aBA/MFC6KdsdMq6ZqfT2de7u4VgcWXgty1wNmFiTujnKd3As65q9Xwhlpof7QxCLKKbCkg+9Q90hYR1wNxZR1VoraEhIewD4S5SH2TxQhfJwf4x371pdue7LDDH46ZP1gQZyxMwCK/0HL+/dvY1Ola01Ue35vH6Nxk3gyp8bRCqKlUKYzN1ak5SYaV0Xv6IGRYS5CUvOKa+Lu6l0DLTHX7jnencWGxIAImjGSHT9wnDtq4C7D8aUskgQoQWopkS9DAWHECosLN591gp7t7Bcf3gEOcmcC+B6NSFr7NashQfc7X0V6S9zb7U+vnnz8OLl3d3D/cN9BFm/WwYRCYtq6u0YuCd7VHW2jcXcn4RxVWXpSx4zEFWXEgqQ4p2ilMLSxyXNATG+DKjBKv5O7QhOtxNVojd7/fYPX/3Sz7/0v/aBZhV2d+ckSVWTLnkJYhCfY6xX7uFjrRpYlzCPUursJqo5pZxzXlEDwcwqXESJwoKKc07rQWJv9NWFt/azf+O6xS1ucYtb/H86bgL0LW5xi1u8h/HD7371V/7lP/udX/9bx/tjtifSxipukpclrwfujyXCqpKT5EWSDnnIhUlESdkp7Lx5qeQOZoHVXcOilXo+1VbD45izB+2nLYJUE2k6PHxoRf70u3/8ne99+vhUglMwnsZhchwcCYoXLx9+8Ze++fKDl622H3z/h29eP55P57dPb3sjehYonCSszWAXjQgz9Emrz+ctp3Q8Hk+nrVld1hXHnlJa1shB+14jXPOSSYl4r+4WxLztFtHg8YyInKmx1VJfv3nzfHqGiPn/UswaWsjG44l/NPuD0KoseFr+iwL01AiYBeL1/IMw3tglaUhTNFEV/M7zecSFCQC+gYyC7u6C84CLUJhLrcBoJNUkag1ZAFdN06fWOdbu7j7L0mOUKuO/ePATfDI9R8nwlJ9EBL2SoCZDq50iNRG11rZtW5YFHkwiYpaUEpSg8/kswi9evMDbp/kaG4whr+MsXMttUyyY2zQzswaSAwIK+Ox7Nq4oXx/CtSkVrzwcDkQEtVdE0JVRrqgLUBmAv2jNRr15l4m3bV+WPE/CFKCJyMyJYGjtUuOUtuOSSOhaNhGVUnCGYUo9HA6zNyN4pNhUGtLMMNLKdMWmi2oDS+/FMozh5m4Db9BxvaA5M5pneh/MF47w0EP7gCGKwZ/t5tP+0hhKR4x50J3OcB7TONKY+soVBMDdrU0wK43iA6IBusEGeLAN+hzButP1VxaVkWIJSIGtVSZWUYO/s1mXzLsUe2HCwA5cS12WJedso3teB+Ywc2cENfxuoK2PqRQDdhGjDV1KCQUcEHEmrUJVt20josNhRXbhdDrVWnFZmRlCM4Yx0hkAs6Cz4nBNRikVuZ+ZpOGRBMKhTTjAnBEzhcAqxATNl4jWZe1nI5x7jzsnoiQ6Uztj4Kl7lFKJAj7lqbvVWvc9HQ4H7N6k9OScMeDn+jCnHt6I1AsadWI8I9y9NUjSAlB7a829V1oMeyy5WRu9GVV0Paz4CKyWV8pbjKUYaAgTFk2aUjLrWOrWWoTntNCAIGGsIilzkdTvVqRzxuXueRgdFSFY05Yll6IR4In3ucYiquzwCBPXWj0854z0jYoEDSpNV88FNu3Jd8A17oMkLdu+ufnDw8NIAPRRtywLEY9unJc03rwz4fyrYmo4GkgiRTNc8DAyT3ywM7OorgdDuuNSr9JfiT4BPisb0KdWVChGNRXRbH4314hpWhdWEoGV3t11Eq47LMdFkBC/mKnfvW1jb2BhvlSxuFut0hrXQhzR3NxBNaGx1vUGiU9vn9b1mD/I9/f3zez5dK61NjPWhAQc8kPmfqlWools6jeggNNcRJiD0dYCGRqUCDSkWIIoWt1LUdWUQpIGB3G3OmMAk7CohEt0k/ggChExUSV6rvajV08/+eLp6XS+u1ORCC8imlBok7JqitEaGF8J3L35SJOOfyPIWsNSWj20tdbMW7TWWr9BqIoEhQe34Hzkw7q82c6telb+r/6jf+ff/c/+W7rFLW5xi1u8p3EToG9xi1vc4j2Muh1+6x/984d7WjhS7Hf3RzquXltesmoSSe4eTCkvpOrEtVSjEJGwCqZtULi38/OJzJJKWGN3pViVNdytMfO6Lse7B2feSnUS0sTLSsvDq8+/+I3f/t/+7Dvf6x3SJ/+5K6UBPuXHH3/8q7/6q0n1Jz/96fe+931mPh6P5/2MJ+S8rMTi5qIpiJs1dOgSETwe19pURJIeDodqKYLwoEjM215O5w1myefTWaV6xPl0JiJRPW97uDczEVZRNtu3/fnp6fWbN/u2/UznfYhcl1ririVfu5qDrkxkg3gRHMHDsdkfD7v2RkNOvhCfCU+7xN0UPdsPwqPKLB1v+s6D/TuggvGzjG6ESVPXDvetVc3LsqSsqqXsQ5MCS7eHanLv5f8QI/Z9dzcYsiKi1sqdKeFmHuE5Z9U0HLu9RRges1X1imDr8C22VmFwzjlDe8KzPR7OdTQzHCpt13CxS1PDvVycsTMRDXZsSHU6KschJ05BCibWZVkhXsB3n3vHS5sC3RS/eLjVaCALIiLnDC0MRzd6A+q6rrUW1Q5PwMellI7HOzODGgq3spnlnJdl2bY9IqDTmXmtFTTqqcdBoZ7S4dSjp5g+VPKAzIvLOnka7g5X5jSMz7mGkw9Id4TnYSmVoXpPBWfyFkAsxV/MHQ7K2poiDQC8gYcq+sB1VVukw5q7Dq09YTJn0sAR2BSv+ySZ8wWKtvC0Y9Oozr8eDKOX3rBWj9p+6gAHvHdYdjtYIHc6MPIoFvPCQbnWnD2ilhKjAgCZmGBSVRXd983MVSTlTETn04mZU84pZw+vtc1zOK8gNg6ISill+MQFYJCUUq3t4WFflgUm0hcvXlyPRrAmcs61NgzUnHNKCrGIKCY0HKfl4eEB+RoUGbybb+gX2odVvB9+9J597r1hKQ7Bu9tR3Z2FlpQj3M1qbTJg5cx0OHSqgF+1ExyzsnfMg1COUNVSS4TrZPgM9r1qgtG+NQcBhoZhXETXVUspSGSqppTyGM8xdf/dTVXW9TiGLmYTzwVn30tXWg3cbY0Qd3wuDMs6JmMzc4pIOSVNpdaIUEFVANYBUVWws8HzwUxJo3coCkfuH+5wdPf3d0SMWh9m3stOxMLcrAGRdHd/j06w1OfBsKCqunspBStz6TJlz9J5QJxlEbnXuwhvrajqw4t7a42Ij8cVqmLOWJpoWe7cvbU6F8OUMjG5e6JMzGZOQYuswR0upPplagqKJJac6Mp1LtKTSypKROauw5Vs3p3m4eTu6EaI98YgmyMRgvmONKyIuht2G9eoWvOOiu9m5Ojt8zC1RpFRXyXIfGQrqaNFWsu1pJ2oRFA4mmmQeH/9AH8R0fl8fvv27bKs5r5t2/l8DqLloDDoozAC02EI3F09H/d/ju4o73/DwVrPgDn4W1ilLTwiqrXqJpXn+oXMCXq0akrIdJEbcnxQnwF6B4jj0y9e/+n3l7tf+Xo+LOTmpB5qximraDIPEeLEeeDAzM2RLuyrQi+sGgStgswLi7bWaqtmjdklaThTUAoWr8fleMilkJ3zUa3RLW5xi1vc4v2NmwB9i1vc4hbvW/zm//jfvfm83h3jow9fZqpkdEgqoXDasJu4Ex74rAaLUZRtp4hlyW4N3bIivJm17UxMpMnh0xGt4UYUeWXNkg+x3qnmuyMFJ8oLHY6v3+4/+vz5T77zw09/+tqJHDW0RMTeHwwjROThePza1772rW996/Hx7evXr91tWdaUEilBUNOUicQ1SBSGWlj+mEk5HTWth661sWgaeF9VIRSAm4tIELkZnDu2GnM3Nroza282RR7b+fz09LaUDY7OL1cB/z+NUe4aw0PVRc3JqR0/4NWQmuF4ctTycpAHdWlneD6Z3VmEAHCQUVcrzqwk4jwc1tgsttPF7C6HT2m7i9PIAHRMLkOFZDxEEiecREhy41H/StDkGCXrKkrp0hUQhdpTi+QrcK17WDMXVQmFn2s0xwrvRyAssLNNqAgNZQHKBQ0VbFrwUkqt2b7v127N68ArAUSGfABtdL4Sb4QgTkQQd2B5FhEovMxca4UQhhe31pZlYSaI7FMrpCu17gpBHtd/JCKzdjrBotvVXhpUBOhC10rfPK5aCxHDMN5aG6RygpG/pwfocnLA9HB3sw7LnrRoOCzxiVAKJkoYBtJ58rHPQC4QMYgZ3ftmRlcNADH03u2d2Y/aB7PD3JImTRrDMKfDzA6RWC/iS5+IMftkjikWfZN9OF4jSGMMki7D8fVUnJP0y8bofmjY9763F3h7XGzLg5PeEc8kIkzcrFlr7rEeDkRUS+35JqJWW7OWNEXyUCtld/NInTXh7sxkxqJi5rUUZICgzjsD2OLuUfcSFFidmHk4470BaJsT+qxi7rNw84bDBK6gWQvq7CMPM+/Xymd7UiKUzKt2Ykb3OI/OgYy56b1xY0SgcSLSX8QX0ol7L8r3cGEJFjcjJ4Oa1pMrHV4cAQL4pYOoiDSzmXKIIDdXVU0a5tVLJYL43q4YKhAQKQJokE4IwWl0SHXMJGY94zVWJzb3iChlw7BpZlgsRSyCRk2GwPIsIq02oghXcwsP5i7chzPY08OhTGajSWlYZcxQiuBoHcWAuoRaG6Tqvk6GWzPUi2AgWlNiDo+UNHrOLIvwvu/dPm+G9F5KXQ6mYcPnvsR11AkSfhFBNFcttGbtHe0mRUFEpJROn1d1xxVhM4+gWjsRHnzw6/WNeylAMDGLYNrD5CsiszgG0xOJPWRjhwCNwoiohL4OkZKKCEUAU8NsERSGPn7svSFo70fZ7xoRROQ9LcLuEw2hqt66YDrqdWb7BGR4nfSqmud6VeEhlEO1v3oB05gAnWsRRMQRVEp9fj49PJToKPxq7kQSQR7DM2wdpz4F6Jn1wb3G3Dv6mXs3ziYNuyGakGo29yDCMgKKPVLC8L8zEZZv/AeroKvqxBg5kYx18bPXpz/63hcff/hhvFwOVvfznkVA0Ug59yIole5jVuZRVyICyhaJimq/jY66JSbm1iy3ZN5QLhCOpVRJOPLy4cP9q+ez1X0nvbUivMUtbnGL9zhuAvQtbnGLW7xvEVxrzcsxvvJw79ubyiwUQsHk0byzMM3cvbkD8ly2TZjTesDzCCQoDc9k1JHFyiqSczNjorSuko+Ujk1yXg7Hw4EkU17oeP+9z7/zyY8+//6nr1+/PcdQWPt+McECrZI++ujDr339a7/wtW/86NPfffP4eHd3UE2impbUOpqAPZiFWJiCmclhp/ZQzcu6ouVarTVlMmsyPJtTsMPDpxlIlLwsCaouXG8RUUtttYV72fftdPbWCIoW0V9eg57GZ57yU7dU9a70Vy+FhIMnN7ixoG4ROVkvqB4a9KyHxyFN7dRZXRSGLeLRPqvvQgzCYzdBz8/ngZ2eIhaPhoF1EB4AWm21tVJhoBORcG+twbeFZ2SHrMNsreG5WVVUBYgJGmKxdXWzlr2gQdiwZ3Z3ZC1VVUOkefXRPM7dSrmwUODbrbXNBmjwIUIHOZ/PYB1M0C20YHwys6jCNWzQi689v9haKQVcDqJsZtu2gTo9Kain01lV13XBr9u2YaSdTqd1XZdlQXPCiOidplqjoYTqaJ8IRxgMa+CKoB3ikH0usq+IqgpAATD+Y6jDdQ6xeCI4Sik4Xnw0TGdy6bXYSdnrem6tTZc03JT4JJyZfd/nLrXWzGwaUQHCdo+cdZ52rCPCDET7LHIATTWmEkOQroDApklZcXez0DRIDuhGqL0evRcLBLzKBBFqLCXcQRRDDgYfnYi6tETz/8aEfHee9kwLETHJxd57JZ8PQTr6SzGT4bikKXLBO19braVYs8PxDpqRjIqEWqubr+siwkGx7zsF5WV5ZzVgTvuC7prrsgB2YaNLIQ/dlpgkvQOodfdt35a8HI/Hbdu6wXldRWXfd6iBsE4j00DT0suirLDDwyYMHgURqcpkziRVFa21MlHOubaObcF20FORmPK6cLfBJsjHHMREk/GCedGSXIt6zGytUhCzQLcqpSDfUwoAzZHzwsStWUopPDWqrbVmDaUPHfjOPGnyXzqrVXhg6qEzB5aClJKZQZuTJMR0Pl8o6twP0AGRSJqSavg/43aAWdCVvvBSa6n1eDzOjA5N0o7ZsiwqEhGltNbwX0tKad93VISgyIBGPumw5JnEGofJ6OeJ81xKoc726edVBuBongEaSS9mznkBFH5ZFszuWZNh1rN0pZQIPx6PWBCmj34e7/UGRfpSPy/x6FR5ARbNd9G1omoGA3heEqzfkPgjYjY1bGY+yghEhum+b5DCe6GJmbEKX90bx1x2or4Q9N0gEmbB2oWlZPzfxZoNzHRn93ePNn6d0Hu80VtrpVqzvmYHUXBc1TYham2n0/l8PqeUKbg1r7UKiagGUanIVAk6+zGj+sLc8E1JRMPdrVlEsAihK4B5Yya3iFARsgt1hNHAwCyISEOEHIinjkBhUWHpHQoZd9qZj+NeA/LTx/LH8fYbX38SP34oJbZnCV+WFd8EjncHTcLCklNKoipLV6EJAnVE5GXBCh8RqsyMN7BnN+skH3w3E2ZNOTwqywcPD0+lnZqdqou+U7p0i1vc4ha3eJ/iJkDf4ha3uMV7FX/wa79WitmhUazbdranN9ubNxuTEgmRRH/KifFoTnAUq1IQPGisojmp6CJ8EGZVVmVNoiqq3iyI03LgdGBdKUSISQc5t8Uf/uG3/5d/8tuPT8/9uQy7xZ0ZIUIelJb04ccfHu+Pz+fTjz778edffHE83JnbXms4wRLGIhTsEWmIdAFvnYc7oZKaiFAKDQfc/AERV9KVhVPXWTx6FyANjVbq09u359Op1dqf9P8K/uerit1e+3vZBKpmh/3ZCe2i8LTcwRYD0EGMVw9trEvQQ8/Gr30XWViFdRpD+fI6+LH6uR/6xfyELmyL9FZUNEVD7hJeQrd6a4FK6iWziHvYkBticFchMJk7hLuUEhOVemmJ1prVWgjFw71zl0478/TqIh0SgwU8ZRcdL576A/Z+SiEz5XA6nQeag6Hw0lBkiFh7vzIy673XoMNS1xC51oah8ubNG+806gTzHRTAIWR3lHNEnM9nHMW2bXgNnqsfHx+hxcAvDMEopQS3m5mt6yHCT6cTONFdYbziD2D7AGUwM8REd4ez8s2b19hnHCNdmXtPp9PU40BHwa/M7G5ffFEHagD2zFjXlZnAxiXilHTf923b/Apd0vWgITC1xszRWoMjMufcwk/nbeZF3tWdZYpAM1MCbKuMxExsF943JN9piUVyACX4l66aA1oTV7+OSYT5BnkY5v6hBl10ZR5CdjdH85S2x35fzeD+QoiMw3QdqsoDbh4Uvfea+/PzM7N0J2n4VOQh/MG6TcS1fanGnEV2jLrWyzh0Hv7lEjM5v7MyRUSFnOlW9oLx0MxEudaGZnHw/F5PKKQKmLqOvO/73Bp1dsSVAM0COscUGVHFj1lgER7erAVRrXVZFlUttapI1jRt9YfDgZmfns8ThBJD302qy7Li7M0SFnhyITsScSktqcoQHA3OayYZPvToxRRfrn64PlV9WnlXoK11yrkkQWLAhuQNHgVuK0CBMzNWwuvAegnrMRGllD28tfb0/Ixedt691QV3h33fpVcb9FKJ1irNDoEjZTUvRCv71XUO98g5EfHsU+duTEqjaSrNuoG/EKp9KUaW63zecdtpzamD2tnNT+UZa+nzc/9h30v3YvexoUizqQruv1hAzufzWCeGPdjD3WprS84Y/7PQBEt6a1ZqhZubmMu+wZoNVo+I9MVUeNs39+6VZZGkCgEa8nRO2lrtc/DqZgcsNfoW5pHxwj7OkzXkZFIV7WumN+vdNceiOss3aEImOpijVbeeyJ8y95zRc9y52fPz88PDi5cvXxIT+CfYTF46nApFUj2DBjwJ0UyU9hIZZlaJnLFeWDO0tyWi2WiUmUk4iADkICJlQS8HH4M53L3p7mZxlZemrtkb0R70tvoPv3j71fv08x+/CI7ktq4HZWYGQ6cFeRQs196R5O45J4Ct8rKsh3VmOpMuy7Ie7+5SSkkXVUUNVxBFL6Mh8uAgUeHa8mpRhW5xi1vc4hbvadwE6Fvc4ha3eK/CH2R57fvPVfHl6Yuf+PmV7adGlFiTqrASkcEMo4mJCKXFTJBOJQGPuWpKv6LbGgAAIABJREFUosrCTuHheV1VleELIhZNEeLevLZqrVoLSiX0bdU/+P3//ff+1//j+XQOeueZHTX1eEg+HJZf/OVfvH/x8Omnn33+6tWbt88suUswaGMUsSyrh5dSkzsFlVJZhNE83ayW2lqloNYqHsByUjAPxvNjx6TCTkrcK+XxbNaV09bKvj+9fbvvW/fT0aj8/6sENCuG/ju8WDxoAkTMwcHMMZEcPE4Mo/kgOQ2l4+r/+gkc+zf+W5jkqova+LfrgNhe94RCaOPuchp69BBysdswn6JXlbA4BUVwUEoK9c1hkYaEdGnEJx5GzKqpl9KXKiopJWJute373q/HYBl86awJMLKQ9pKyCHgXzJRzRu3/dL/OJ20zb9ZEJGla12Xf9lJLb2LHbB1nka9gx8LMQBb08vYI6Fw0fGvMDNN4eIzGU514MjUF6E3SVXJKSTFgwkNURLSUPQaE1z1qLdPjCdvvumwBQUpAXJig2+7gg1TdzIC87XhPimHHNijj0HqIohdoww9InFICj7WUykwqKqqolwdhgzofIOC1NGseATCxmXkv4RcACqhDF4hFUjNmcjfgF1QUFd+lX+Kp81GMBnQ4Y+bIaoxSend03WSwjGnYkHEap06ECzRaGGKoXiQT+PbiYnLmnkEJFMQHdz15Wh15wmiurNS46FdTvqvWEWMLUMKYe+H9YHMz9Yr4lBJUazcHygB/Zw5kPlprQc4D8GL+JX/fWB8iDK320PsRwBYIx7im8U5/1IhorWnVVlurbciajUXMLdCYrnSww1TDe02K9/KMzjtS9dF6EQJ0pykTQyFSETTMRDtEd2MRB1OlKRFVMzMTldaaijRJ5mat1dpQV7HtW8TFlotsIYaQDRWPh88XmjK079ZielRhZ0YLuwmbhov2SwsLRO3RIbIvO625iKaU3DqHQVSIqdYKdba1JqIs3IBsHjOLnOhdkVEGcdjMiGJZVmKGHkno2TgGcEdDuBOzqrhhMknnL/TVWGYBBMZ7mEkf+oyjbi0hl4B1z92ZjZtfZxc6AuUyrnDRNaKjfsZpERGhKIODzB5Ra8k5MfdmgympeQCtMNZebq2ZewoFSQNdMa01HOPQ0JEds9ZHL5vZzJmhHAR9bUFhIeogIyz1EKCBZBZhsMtxwkXZRKlT4IOZwxPWE+bLNKerpcBao5x9gPJH/imgfmKzztwu1umI/tHCYxSNvyJtEihgoiG0A6ZMY4l6ZxBSmNvp+XlZ1oeXL9d1ZUC6e36s86ZkloaxgL003dwzWQuQV4gQEZIxbCQiQcTkaA7sHcSENdjDg3tvaaGRXiImcmFVdgsK8stuB5ET1aDnZj969fjXPjzG1z9c+X7lOCwLSujcLThIwgHzMdPo60sz83Azq61t++7Dw64pLXnd9rIsS0pLSr3h5wReu0cNejZtpVptUhPl9l/+x//Wv/ef/kO6xS1ucYtbvHdxE6BvcYtb3OL9iV//9V9r55AX6aiirX3+4z/PvB1WiZBIyimTqDObheZFliXnhUkC1aOqkrIk1ZxTWiRlFqWwsp3qdkrHF8wcz8+cs4hQLe38tJ+ey/m5bWevW/D6+hzf/vHT7/7W7/7xH323ur+j446fzEgT3T0c/sW/9TfX5fgnf/Lt12+ezufi9gYiS6kNBM9lPbrZ+XzmTSANoBUbi7RaB47AS9nNPKX08HCPwmEiwlPuxYJ3PGpKpRZvhi5YkO3c/Xw+Pz0/11qI4Ar8v7HR/V9HzOdPHsrY9bFfynIBG+g/0XRzEpS0y1PstZftSnIbW4VcJeNVPGm2c2M0vNwx6mu5O6DB5B4C3JVsM5Xl4QsDUUO280bjodfda9khN08YsUdo0sPhWGu11qKLBeI+pD641QZ4gTzADAHEs7W25ISC3giyZrW24QhmZkbnOsiQ5u4eOUFScTNvzVqr+763WtOyDtBzqGoyT6pEUUqFk7HVip1Pqu52Pm/MrCopZ1SGwy9MEIxG2TjLgKYQpaQUUeuViZWZAkIzq6beUm/Y7FD+TzCfRpjZW4cUIpoSnIwXD3rvboej9K4A1sqClE8ws6iWWrF70cu/eeh6nSwqnSTA4e5uMrosllKvzcDn8/m6zHzmKgTqMDNEJmt1OR41Jaic0/HHzHBTRkT4YAWIMLM1m6pfREQ4czfCX41GJmK/gvTwu4P8SvgfyZKrcv6rJMs706RPK+kM8Xe2OVNBlyoJGqmH8fsUSanXxXc9ehiYo6vxrP1CU+Ha52CH7oY1J6acFWX1aONJROu6cPdHv+tl9j7SsHzlnLnLZwCFsyZl7hfoOtwas+yyx7goWpVFsJ+4AB7h4SoYt1VUhcWbIzNXSyEizQni/rUDumu+0bN63oDm7+Ijp+77VmVVYeG9NEhOQlQGl5aJTueTMBOTmUOfVRFVMXc4YeFHRkc7IjJgcXt+i2FCHlcSo+lagL5wKt45pYMUwcKqihEOKy5uDbgioso6pMaIbduZiFW7AJ0UI1X+mfeFDqIxqJEs4hSt1iDSlAbLu6tsSRNRbJububAcDkdQdMyaqKomawCPkKbMTF6rCGuC3uo++rlFDJhyRBC7Q3Ee8iIxMqk00mlEwawRHcg7fOVE3XMdIv2NuMkGRWuT4bMQsZuzCFFYa6IqoqVU5Km3bSeipJmCzOx8OqWEjpp9H/ZSL7UKxLVWounxp9Zs35E4CcE9Zel5u1YHLEikj2Ezb9GoYpBgqbRWIem2weKn8eLDYe2DGa+rLa5Y1bjcIrz2vrU9DZOS1tp80KiJaFDLu2Z9KUoYeS6K3mjhagxefnJvp9PzejiYVeagiFoqcoRIVRIxEl1zDEd4SkzEpVaKjuMIJyd3d4rQ6BxtHwcC/f16IuCfJEJEdfj9IwIZQFFxV6xnX9rvRnRu9tmrN59/fF8oPnjx8CLrKiTkgpqhrCkrKTm5mZOFN0Mu093LXkotpVQ393BzI2aiZ/7ibUoppSwq1InkNaX04sXLWuu5tXOlur5oYbL8n+y9S7MkSXYe9p1z3CMy761390w/ptHAPADSTDBIa0kLSsaNfgC5ljbgitxq27+BXAEbyrihbLCXTGYykWY0SqAwBgzBGRCawfT7UdVV3VV1H5kZ4X7O0eJEROa9N2/V7erqR/XE1zPdeSPDPTz8ERn++effcWs86R5fnRkzZsyY8R3ATEDPmDFjxncHraXNsh4Uv3PnVutdqteEmiaTQHJumqZ14eroi+W2zU1LEDN3c2kaFo5ZbCi5au+Au2rtN7XrVp9XUtXNOjUNM/frdelWtd+QV9Teak8pPXp8/Jd/9cuPP7kX1MNFFXGwPbfv3HrzzR/cvn3r6PHpRx9/otVybomG+DkWthDmq9WaiNp2gcHXMuwgmZmVCAhlbgrRFhGnJCmltm0nyVLTNJPai4UP8oGWWktt2yAx7OTkpNtsdPATYB630j+tmreE8nRb+z7v4SzcL5uouo9RAjE6aAxnDGSyD+mHo0HADbrps3U9BJ/yibejYNXOlcfHc0Z7g6kcIABVTanyWFyKDePupkrE8GqT+QncVF0tIjQhGEzhwRd4JHONeQqyxGEzPTZVp7WPbbk0xMtydwKsFAS/MMrFo5a0EMYYigRUQijzte8Gco8ooh4qhZpQw73EzEHsrErkZq4Kghq5lvAjMapETMwTo8rMIHIPZTopY9TfDSYGNNIPDq/aB1M/8RQ+ymsn3etADLlbKTaQrEREtuPMEG0R6mCPSFs+kAimipHB3OV8AbiFJ6mb13G/edDSNcbIWZUluVV3B7HxYL0a7jyuFnma6hC/q0TsLh3Vg2PHGXWC226lNvS7871tkPYTyGns7YCPW92jP24J5YuPj50vaBgnO9ixznACiMewYtieSdvMaWcAbAlo32Y+NPqYKLKxcU3HiHQ7bqYsaEtRA6ZB95uaRnV0mw14JMEnXjxGCWhUR7rVOg3dUMjW2u+tlGklYGqCWoho0IVjXBBz9zru8KdSo3kGzamqA+GuE8sbQ2i0SfyL0QMihkMZfUBq1C+0DK5CYcRDQ42Rh4vuZA5EmFZxhhCBTlNPJkLX2cQwn3mMEmO3ysYHVpD10+2f5/TjSQWEc+6wimBKNNgQDytMzMSjKjYyIRDLMMq0DlpU9/N1H20fLUvUbTaDuDyM/SfT7WDhmSDm7kG1G/E6lphia4NVq3WqYQ+ffatGFHYj4cBirtEliJh0GN1ucQkHYKOR8U61AHCCevDLbjQuzMDhVh1wJ1ONu9NQe7vGtoWiA3c8qMAHI6AKhxKYaGB3qSK4VfdaS0jUhxFkGumjg7k6CMYcKuDh+eYI4bZb71qGdSk1j1swjeB/U50PQzzCa46jbwiPucMv911HIR4PY4rRxXu8fXeYEnVq7oOPilXWwuGrM70EbE8fN3fsHp4+7cf4nKylOz05Ykkpp7gLNY81x7C08jE+LYBYwCXinHM4oo0bz6gvxcyYSHKmYTnWeNiEMdw4jUFxp8+TIzNF7F/icF7WqkOY1p09IPGqcbTxu49W7999cO3NV68fZNXeTBmeRSS2NwkiRqYkRoOmDqF0QwRQa02SYv+cqqo6nCbjtyjbGEbSYtNR1UIomaHwpjRNrv/mrX/w3731by+v3BkzZsyY8UJiJqBnzJgx47uDJNTWRVrQ4UHbumm55tYLeyJJSVLOLsIgSpaaVlJ2g6s5wEwEVy3QgV8bZjO11r4vfderea1aS86ZmLrN2qzCK0zJTVh6w4NHR3/9y199ev+zQcx7fmIWDKN/73sv//D3fq9tms3ms+OjY+a0bBcgqLm6sQ8bVM00SVosFkHhiAwh14jgngGE5eiQ88jj8U6Yo7AhFpGY6jVNYywybhbuuq7v+3C8dccof37CbPKLwndnyOePutPZgyPDMXFkF3jt80cmOeeZQxjEWDTJn+OLsxfcvcygALVRThvfR1rdcoJbvizEmEGejJe2XivGHJyNjIc5PxHcPDb7hkMvCGwgUavBMtSR19zeFABgx3FguvcwKjnrtO1BwkLV4GEXSk7Qkacd+YSgA9h1S9g54ORWgzaN6TiDCTayEsSEgYsESDF8mMR0wRAx8xCwbqCGd5YxiKYcJrPiSVUXxGXQ9OcJZR8oOxo2fwMAmQ4a9W097bAw0fLhm0E8DLpwACXb4X0BgptGJwlJITHHjnJzkNmwnd8dINMKhQ0UCW1vjAch9q7eGQ4a/Hlt4tfjXgYTcsfWNnWy5tlt4qnr7uDimg/tstDuOwT0xIAPA2ssxpTpmYGzc3z36xi8PlUYhm0Ku+Nqt1SEMXLhYG9tFt4NY2ZeNJjmrcPptEVhLJIDCFcHDL0l6FHDhQo5Wx9nl5cuLn6NHRXnrohoX0V0PBuWGeycKflIa2osZoF8fHKY25avo9FlCbRD4o3rBVs5+cCbR+ZMDCILsnLk7Hb2gOiW/yUgXM7dR8F+DL3zROBAmsf9TWuKZoMCfdKKBhU+LJiOzyuyuKKrE49NeY5opLG9iIio+mCWQhzrT4rRDCEuUs0RjhCxNlFtrJNYjdnm70Of2Y6I8J5y1XFoGYyIGI5JmwtgCKw5LX1Nnjhj9zC3nVpFNNC0KjAdnbpL8MtDmwLTUuL2xwoASL2ChiZ2wAbHc4AIAwHN42CiIJudomls3JRAw+6NOvau4anJHmYP2w4WRbMxVvDYGAMDvu1xWmyqzW3Xm0bu+HNTo63H7hV2y/HIHLPmMQl2G+US5vnCwBvMZPqT4+Nr129E8ORSivUlIiJMMRV208Syh0zxgUtRMxCEmcaoicOSIbO7C7MD8e+wGrcxT2YW5rpjmQUGORErIryzO43VGqU3YFVx/2jz3iefvf69l68fAJtOtAiszTnqSwYmnZkTE1k4vAmHMYeZNW0rIiBojQOmqrVqxDt1+Bg7EaoiSZwZC0FuNsoKvLrsT2cn6BkzZsz4LmImoGfMmDHjO4Jf//n/5lBa+q2bd5okKGtKS61k2hu0au1LJzlLbpomu1ftK4hhDtP+9LSWvvRrCapMq4BC4lS60nU9HAQmllL7cEBs2kVKh48eP2KS5uDag4en7997/Ldvf/zZ4xMfeVACxm3pIQ4EOV579dXf/8lP1qerk+PjJqec2pSyiDhgcFOLydVmsyFC07TMbG59VzgxM9dam6Yh4pD5hOLGHVM8t5ie5bAKAXLOfSkxn2SR5DDTUsrJycnpyclmvTGzgS0zvTL/vEsW79LWF9PvIbWnuSxtj5z7Zpv47EV9dMH1YErOZb0zVT573XE2PeV5hu0b6Lsdqm2b3HdTDKxVkIznyrrzyYO9PZNT8FLO4wlKNpDiE1My3iOeBB8ZxbN8k7lvWUfdYdt3TxtUi+eTb4nEKKjCdnTqbqMrw25twLe0hcMRvSioi/PX3VKjuxzJeFX3cXBMauAz5Z+uvC0CzvBIMJvKesYKNQimkXeJCjpbXeNfqkRx1+MVR7+J8YTdm9ppaZs4RdrhY0bmeSsXHNi6HQLMMfTe8flwrjtdgjNU2dmG21ZZ7AzYKa3jrEfseCSufJFJ2mXptp/GPHbZ620lYRpeoxo3htSOVjI++AUnjX1PiYnN333UXFY9F2mvS845W9ZzaYcFjHEFxXc72W677TLwZ4o3tsP5x9t4+2fXFabPRrZTtrF29/J7HiXT6Xw/O1rO3PBumYf/kpv7SBZHJhPTuO/S5NvNPBcexhhu1ndKPlK0gxEvjfr5MNAH88DD+viop52sLtzBcClzd6VgeccR5dCdrjs27u442H413oJvHye7lXL5U9eHbMe6uvDLQpd+5Rh4fADj9pHxTPKhxacq3B0g8Rvn7uSkO8XzbZLz48XPd5YLf/pUdWcTnl/WvZjTWeP1HVB0qLOVcTb1ePd9v1HT5XKZDw/bxcHJyUmpJeUcTLKNDjzRW8JExUf76cjJzKopM+chum81s7ZtmQbvlLANoZGYlh0XkWkVBEASAbhqAYOZTRVwHj2mPBy6HAI8Pt28e9d++OaqFdGjzxuvDXmbU845N83y+mHTNJIErrFcCyIhhgMRIDkW4Ry5aRrAapUkKUlE+BhWhneNRIiVxCQ/XK0enpb765Rl77CeMWPGjBkvNmYCesaMGTO+I1Crwkncl0nqeqVlHTyss1u/MasU2iozrb0adGQb3J3cXatqMVdyY4d6+C0AVcXBkokFICPjxO3BYW5bYeGmpdTmg+sPPvxP7939/MHRZlXU6cwUflBYEtpFe+vWrTfeeOPWrdt/88v//N57H242a83I5iJi2/jvIVJWM+02/eBGSiibYqOMNOwyAqH0mbZ2AoPJ7CTMLLWqWakF5mFA3Pf9er0uffGBfQZwYdb6dPg+1uDcCRhny3soUT8/Zd/Nc3deO02dz9BGZxPuvfSeg35WBRe5DQLl81eczDzOJJim8pezYjvT8vEDwWnvCTusyZVb4OKJfqGYXyj5ue8vsBA7JPT+TLZy5n1le8qln5zkqdipyj203YWWiM9nqyvo5t173KeL3HfpEFieHwd7GKCJzaLp0Jm+fZ45Oze4LpRgd7z4vhN2j03C2j1fnU1CuFA7O2soe7I9W9ixVOdL84UfLt8MzpD0fr5d95LCz/eiz3D+dug9OdEOkfp1wacxtbvn4swZe9NdeIzsu8dz+yCuWKJ9Ry4r097M9548Pb/P9p/9Cc+Ojj01cHEQnT9p7wLjE/HcG923K2iXtcPYjKH43WzWTdOknKMZN+uNI2LPbpli91Gx7uHAX7uucx8U8jqG1rBRwh/vObVUH6PR7hkI7lUVDhbWYNkt9jsRORDuSMNyzvCOYfCT3j9+XO897u5cO7jeHrKuyaqB+qq9bnp3SbGabARE6EimsDsTEWlDAQ2kJMIEIBurspoOO4YowtDKQHwDiUBZXJarrqz7pdX+p//zP/zHcyjCGTNmzPhuYSagZ8yYMeO7AP/pT9/f1NO2iixJu259XMtpXjZJGCR9p1AlkHvR2qt5NVfzokGscRIWZuZGtYcjsZB77HPlnJvMuV0Qi6oaWWry9Tt3hBmG5fXb3hzU5vDuoz9/96P7JxsrexjUmKfRtcOD3/+DH7/xxg9ybn7z9tsffXSXkKpSqcosY7i2UaVLVGstfc8iOaembbq+r7WICLMAFJ6Jg8EzU601nDcQAfREaq3unlJSt3BLdFWYi8hms1mv16r14ux7L4P4JRvnomJrz6d93156yp6vnswanEk1knETbXfxinuEeXvLcUXimK5QrC/IQX/d2MftPss532Y8c/mfmPA87Xs5mX2us8XKxMTsnvvzTJ6X5Hfu7126+PzugXOppkW0cSSM+s2t6HOkyZ5Avjt9JU+Urw0vTn/+1g69CwV7dl3nc8xqynLPw38aGf7US+ymvQon/Dzb6Itz0M8Rfub5cUklTfEVwgZ9vV6JSLNYxB6IzWajriLS5BzBb0ut56xv4pVGRFiYI4pvqAbCcLnvh9NqBSjlPTVBABHVUgFkyoNtNMNteAb6qDnHtibJgFX1ByvcfbR6/aVr33v5euqZ60aI1ExNtS/eWa1Va0/uScSHWLsRhzK3TSspAZ5ShDOmJCzCZkocYugBsVugqhITu7e8yDCosWjV/BzaasaMGTNmfJswE9AzZsyY8V3A59f5zQf1b16nLNicPCJdZaoo6mTwSlpglUARjMjUa7Virg5wIhGSLM2yOTjsS6mldGZN07ZNyyAmTkzStkTsWsEgIU7sfbFaOOWqdPJ49Xe/+eDX737QqxIzM7T64C4bEd4JYL/10q3/5r/9r1/+3sufff7wZLV25+XBNXOqCjaTlEXQ930tVdXatmHJ7TKpqjnULKUkkoKnjnh34Z/LDCJOiWNDJ4Zw9im2qdZaSQa/jrj9Ukq33mxWK1Nz7N++fTVcRi1dFERdhaHdc/6FZGeuSDjnm7F7wtP0gJcqQM8fvNr0/lvK/sz4KnHFoXPZysXF5L6PzT2zsnJRWrxzlYuU1GUn0+X5XIaLqsyxVH7utC869p8dFyvxIqH4fBPOeAFxtbali4uxV+4Uzl9z9/nmu+vVhtkUIdPNuq5LKVetcGLmxaJRN2ZucsMc0SwQAftC2940TTiMARAWEVEAEQB3UByTY3B/coCfsAmAxggZ7gSQExGTpCEObZDHNLyoxeKbAp3Zh/c/+/4NefOlpQgz5ZxSJiLmZtGKCNy71amVysxa1UyZWVVLX7VaeIOkxCBo7ReLtl0saETOOaecchYRJjK4aVU/rWnZF0WlTg/c+U/++I//yZ/+6XNorxkzZsyY8e3ATEDPmDFjxncBXfbf/CAtEi8yl5PjRIVZrarCwlqZ4KoOkIOIJImQEEmilDm3nJrULtuDA65a1Rxo2kWTGzIjN4GTJHdTqwDIHKWWzaZuumzy8OT07Q8f/OrvPvjk3kMzA8XVfFT/DZzNrZs3fud3fvD3/t7vf/7w0QcffgSSxfKgbRelulmEZhciSgkETsnbJrMIEbquNzcmDrFM6UGwOJWmrZzMIsxAYkYQ0CKeszK7e0qZhM1Mq/Zdv1qt+q7TUkZq/Nnw9RsU0vjviZ5+LnPwL6zQvMCxzczVbyf2kq3PPC6e2ouemvleDvrZsjp38plP36ru/mw1PrurzjiLL8fonl/QmfvXFqFbj9XuUku32SwWB8vFwsz6UsyGoBfuLiLM5D5EjU1hz0EEIhGWlKpqWI0xETETEMEGw+xirwtNsN8yvFwlZlZmmBMzmAFTgkbcyK3lDsXeh+p+7+HpR58+fvj6bUvWovZ9CY8NMKfkTDQElhy3nTEzUNw95waASHU3cyVOIHHwGM3XzWpflDc9ERHHu6ICjlZyys4F0PXpq4lPv66GmjFjxowZXwdmAnrGjBkzXnj8x//jXz3KSvCXltdasdO6NqpGVq24G+A5CZOoGREzpywpc2JJuV2kdiFNY5xcEklOGWDOTUMpOQHrtZXeq7r2pe/X6xXcmDwJb9brbtO3hd5///6/+/O//v9+/dHnD9dguELdOdwJdyamr7/6yh/86IevvfrKBx98+M4777btoklLODMjQu1E9JyUMg+WggS4uVutZmgkSRIQYAZnIU4ixAzAzAAX4TYvJsNNM2+TqFopJbdNzglEfVdOHEePH/d9565AeC/udYZ9Mp48wb769PsJZz75q+dLgn1h94svQzTO+O7iiv35CUTuk51k/MLn6bTn7OCyI6L+Ggjnq4ynPTd4sWTfKnJ8xrPihWvGs1sXvsy2ou8QpqAU8QlEWvX0dHVwcHh4eECE09V603XmDlM3k5SI0hCgz8PRQlJKkoSZSSSrTnk6EBvBGIh4hntdaAaGehvh0FRNSyE4hZEIweBuCjtvbKSOz476jx+c3n3wSA/SoZh1awZE0mK5TFmYIHAGCGiaJueGiFISZrp+/XrOWVU3m05NOXHQ32GMBkBrLX2ttapZWKXnxE2b2pbaZrnY1BOlRb5ffHbhmDFjxozvFGYCesaMGTNeeEhKZdPnw8ww7U7Nek7EHOIUIZF8cCiS3CnnLCkRSbgsD2HTmYThrlTUS69WN7BwFuxPjr3v4UrE7qamMV0AcTgHduv0/vvv//t///9++uAzc7iR+2B8SCQiVM3dnRw/+eGPfvK7P3x499OH9x90m42kRnIiiJubmaoSgYmIh6lVhETLzNQkM8uZQe7ukoWJhCX8SYnZI8ghSIRDNG3mpkqAEiW3zMxEZrYpfbdZnZ4ed/0GFC6vw67/SfmDSymnq+srz6XaxRO25+/96umGzlcuyWW4zLUjZrlPpxKuUoIrlvKF411+6/FsTNNVUj2Zid497alUNT3xzKdm9fWYOD/7MHqGwj3XIInPZdHueRTkxcBzvMHn+FilL1Gu73yTXcSVf5fPnOi1lNOjo1s3bvhyWWsBPKcERFS+HFQsCzEzgL7v4WBmJhCgpY5BCgdWGwCDnAXuruZAVXUfJNUAQhntZjYtiWc8AAAgAElEQVQGOjR3d3MCgZgpIZlrKfHWZUPJ3QFnQmKC+bqr9x4c3Xnz1Rs3rlPZJLLEZHAisBBMySMKtPZ9R0xuZqYnJ+PVQ1jtHPZoPLzkEROzJEkTpW7uVsy965xaNVJ1k968/PN/+j/8s3/xvz+XZpsxY8aMGd84ZgJ6xowZM15suPv7P/+/1kefZXa26mXFZCk3KQtVBjOlnBcHxMkd0jTM4g43dTc3h9WYz4QzdO03WnuDwsxL350coxYmYmESIWFygkEdObeS89F688m9T3/5t795dLxxkHsokCfzDcDRNu31awe/+8bv3Ll5673fvP3Jhx+tTk6XBwQhgpHDzawUonAmjNDqDgcRjAiuTE6uqubmIIAZ7qoaJPdQfncYuwlRTIHMzc3Uq1ZXKlzN1qvT1elJt1nVWkE0zrUQReWxSvcRTs9rjv0EFsz3ihwvOfObx04hrkQtfSsKPePFwzMTxxdP+PJZfUW4bHA8w+aMK17vax6Oey2/L+K35CHx9XPQV8Gz9fzfkia7iCdU1172GQDMrPT9Zr1u29bchJlAtVZ3dbjWqr515Oi7HgCLRGhl1VBG7+R/4QLVqpkzDz7LIYs2MzYbtoupmpmpEcEcg5pAZHy1cozq6ukVbtWVj+8fv/n9VygtF5JassTeayVCzgKvwVz7IAggNwpXatM6uoKQanUnZ2Zm0CA0YBCnNKx+k6uruRORmRHIYUa8cW2eqXlmzJgxY8a3EzMBPWPGjBkvNj5/75dv/lf//bv/z5/dvHFNrDPXnGh5sGiXi1orS6KUq6FWq1VhDvdatZRipomHXZlWipZea6e1uCsLCYHM+vVa4JITDCzSNhmSjaRUaw+ucV7ee3z//sPTe5+d9E4O5h0lsZurKeA3b1z7+3/w49dee8VUf/5XP//Nex8cHZ2oIUl2A4cdYK2xDZNHN8MkYm61VEkszIml1hozMRpMCj1sDbG713XHCbGUYqpREnMzwvFqfXR8XEuBO12yZfXL4TK98+6M8Qma6J19/08no5/sYHBujnqxAE9Qc58zOpj3U894NjzD+LrKkNl7ofMO6Wf7+dVH1reqw//WsnszZnwHQUTEcnK6AvHy2qEI1VI3m1JKdfcay+buprGCbhE60N0HufP4erPX7hmA0/AuFAS0mxERCdOoiXYbNNCjNNmZkHKqpqq2wz5D3U2RgdNN/eDuyY9eX//g5do0DAHDG8mpSctlQ2TMw2XhIKbI38zULCh1VS1lA4BZeGTHtToR5yYTwEy5aSEEIufcUWoUyaoqrgEn+eZbb7311ltvfU2NNGPGjBkzvkrMBPSMGTNmvNjoV4//7t/9mSQ0OaFbSdsu8iJngar2nUtlLd2qq301NU/CRGaupZRaCxGxgESYBmWKiEO4aZIIszQHt4Q5p+RwFm7ajJydJFdP7eGq0i9+/Ze/fvuDalP8Gh84oJgmweF+5+atP/rDP0wpfXzv7nsffnhyeioplb5WdoCI2M36vo8dmpJSBNhJbqbW9b1vXJjbpnUzVY2Y70QAgYlZzcyIuWkbOGLa5vBByiNCgHotalXrarNZb3ozJwBfjH2ms5+vtql5wBPMBC6juq5CgT3BzeMqx6+OK5ohzJjx5fHk5ZDdMXXF/v+ES+wy0V+V1njGjO805h+Fvbjw6+/jnjCzvuu6Jt9IN4lItZZSN5vO3SRnZjFTBEcrwszMrKoWHHQcR/wDu/AOw8wgmBqIiOBOTgg99c5yO4ERRDeBWDilpH0F6tk7IBCZe+d+VPz+yebTo9N0LfcorH1K3LYZXkXA7AQTZmYZPDaEnSk5exIHDGamU8aDB7Sombl2AKqilA2IweKUOufeJFHq2Ao3n9/4+zc2nz7f5pkxY8aMGd8UZgJ6xowZM15g/Oxnf/L40bsCSW3Dbm5KTLltvZbad6XfhONed3xa+wIH5eTC7uRVXc2JSBpOIpIlJQiZG5i5WUpuJGUhZhFhNjciCJMLGQEVlZePjtf/8W/f+fW7H/rWQnIkZwmAk6Ntmpfu3Pn9H/2k69d3P73/+PjEHO1i4SQGMhAzOxFSclUARkQixOws5nCWWqsZkpNDjGBBPTMTwUBGUAc5kiQQ3ELiY+4ukokIZkakZl2xrtS+FDiG8n6FRNMzuEXPmPFdwlfR8/1qyz/P5Ir8Bai0i5z1jBm/tZgHwjnsXXseFugdXmspfQGcaBQmu6tauxDJqVZiGczBmFmYq6qZT5lM8ud4z9m9MIuASMWGP8lAYJFwjsaY2NwN5AAzCUuSVPZIqglgg/aOlePB8frew+ObzXW1zrvTNifVDK85k7A7rEk55ywiEGGW0AgQEcLBenzfmmIo1hEA3FGqupmrq6uC3KS5frPvXcXfePzLTXv9+bXOjBkzZsz4JjET0DNmzJjxAmPh7Ulz8jLfOjxYkpdSO68b7da1dGqVmEARTXCI9KIetDCl3KRWSDJJQ5KYKQs3+bq7gZiahlJDIohpChETuanWrqzWfSnV+PH65DcffvaLv337g0/uD9OdHU7XHA4k5pfu3H71ey/fvHHj7fcePDo6vnn7TlGTlNvFYXVs+pqbhoR9ZI0RsRGZY6ZiZm5gsAjrIHYG86CvhsPcS1/UlJKklESEKHwPNefs8NL36Dsj8r43hOoHGGQ4z5cj+0K82BXtns/geURDu+jRMWPGF8VVzJSvntVeXLSOOXf+ky+x97Qni6avYsSMp9m4Xzx/xowZMwAABCIy91LLyclpu1gwy3J5QMSl9MuDpaTUdx0RgdjNiImZG3MARDIJmS9zD7PBCIPi3YkymJlEXHV6uQJQazUxIDOcR1H1toxE8XLko+F0Ae4fHd/9PP/41dtgjSDPpcca6paSwGHkThGTA4jdbKG8Dt49vK1FRCSxCBOpqsOZeDQMYVUv1bpSO9WNww+yM04qZFEbf/TTt/7RP37rz77a1pkxY8aMGV89ZgJ6xowZM15U/OxnfwL1W3RjkTir9uvPtTs17SvQdZ3BD64dmHpf1ShR00rKoWsGE7EQC3FiFmYhhggnIai6GzEB7qaDPWGpLAw4mR49erheb7i99s4nj372i3fe/+TB0bobd5cSOTAKXQCw8GuvfP+NH7x++9bN1X9ePfjsMzUXFuEUZDWzEDGcTI1C1GwKg09zGIR7IdNwaiiGHO7Mg7OhA6gEIgKFpChiECL2moLcUKtu1l3pFU5n9qJ+5XTR8yCNZ8z4duFr4Fh3ed5vltL9VrlCz5gx4wWBY+tMtnvUoaWcnp4S0cHyYLlcMNN6DSYGwMzTa1QEEgTDHW5joL/xtSXeeIbtZsE4E01XC8IXQHiU8VY37SklM3N3cmMiZpaURap62XnSOY2vLxU4WnWfH603VW8cNAf5ZsvI5EzWZEmJSYiJQBTb0ZjJbYhryCBmEMV7ppAwiAwgER7e7oiJJUmYXx+YdqprrdpIWrT2aFXc20Xq+6+0qWbMmDFjxteEmYCeMWPGjBcVqaRN7g82aXGjpXKyPvqMoHA3eF/6MPezCK+emtweNAfXUm4kZRICeIiIQ2ACMwFe3WAOVS99cMHrk6P1atVtOhFJwiLp0af3Tk/Xy5vff+ftd3/2lz+///lRr3AGOcidQFtyl6jJ+fUfvPb6668dHCxPTk4fPPhM1ZumZfbNujOQM1eHmfd9zyJEpKZMzMxqBYAwIyZILOFv6OZqZmY550QxsYo5npsZSh13dyoBzKxV+75s1t3qdF36AuwS0NPO2C+EJxDKe3XNTzCuvZj8SWz12e+e6oH7LCLrGTO+IVx0Yf6SzO9zZI3PseGXDfAZM2bMmEDnHxWDhJm06nq1anNDy4NF2xJRrXWIYBF7weLMwW2M3L1WNTPAmWXIncIUmgGYmaqCCURDrOYxDmGtNaU0hP5TNTMRCWvpOMhMKTWW1bTCnYjgsfzv8bBT4LTTR6f98Wbzys0bNw+WLXnyCiuSWHJKOatWVTWDCTGJwc1t8K0GMzFIQGxOsd1NWIjIFCIU7LUk4oaI08K0qVQYi7TsVR+t+tNTlLycQxHOmDFjxncAMwE9Y8aMGS8q2HmxXvRunNhLp65ZKKXEkheH11lS2zYteOFsKUuzaBZLEDsRgL4vpRQmgqlZ1VpLX7q+81qgla0SAaab9crchAeVTBaV1C6vNdK0j45O3//gk/W6mxyVh7h/AUK7aG7fufnmm28cHi7ffuftu3fvnRyftotlKVpr56DqUAezOKBV1dTNiDnnnCSV2pkZiFiGf5gIFAHW3dxrrSIizF3XVdXJGJFomPV1m87caqmnq9PVelW1mpubXazJL4jLiN1zgs1doorOnvDUzK+OyyIEPpl3nsp2jk17cii22WFgxjns7X7PHA8Ql/z5bLisuz4br31RkT272cyYMeNZ4IBV7fu+67prNxbJzMyKqrkLM0L7TKyqfSkACBSbt8wdXgcG2TSEzE1uQFRquK5R7P9y91IrMzNRrXVgvgEAFnBnNyJiJRAkZZbsqu4KULDPU2mL46gv73/64HpLB+mmQpfii5SJASIn4pRJEhFSyjln1lFkTeTwYl774T1NkuSclS1e2cSc1ZU9N5QTmVYwLdumkdYX15rmoPvwXt/3Hzf/Re4/+EYaa8aMGTNmPEfMBPSMGTNmvJBw9/d+8X+uH33KDbuDmJrlQZNYRFiypMwicBeWzMnATu79pi9FzQjo+76UAoebulU1q6V2fQ93imkJ4PAKTrnJbQsnJmJOh+21onS00YdH63ufPuz6si0TkYdihgDg+rXD119/9ZVXvk9Mv3n7N5vNZrk8WCwP3MnMSRK7V3UWIZCJlFrMLIk0uUk5Sw81NXceAQLcbHAtZIldpQ5mbohzTmYWd0dMTGzuqjBC33Xr1Uq1uhlGUc9QjXvr9kot8GS18kX2effz3oR7mbIvWYzLkux+oC/CLM/s84xdTJ3Hn9i3n5rJV4S9Oc99+CJmm5EZM75GuKtZ3/ebzebg2rUw0nBTB4g53DZE2I0wGjFPv9aj0TPcBkI6zDcmOw4mstEq2s0oJVU1H4zLmDk2gXF4PxPcnYlFJKVc3V11d2dYPNArcNKVdz95dHPR3ly0C+8XVBcMTiQ5pSZHzkSUszcKCxm3DcoEc1dTDUq6V+ZwdYOqwZ0AYRJ2ESeCZGnaXLCihcnBDQHU7fDk/zZ6+etuphkzZsyY8bwxE9AzZsyY8ULi0w//0+/+4T/81V/8r9eu3zJYbpY32kYIIDInFiFCLYVJhJlq7deb9WZ1fHxcSp84wvRZhCAnIkkJzA2IJRElJjYALIumaRbLdrF0MzgAbpeHm94+efvDz4+6R49Pq45CmZgS0UhCEW7fvvnjH/3enZdud5v13739dyml1157nSX3pZSqqWncqVaNsIHhmxEEdM5ZUiq11lqqatxvzJqGsIQOIkpJ4mBrjYgcHi5VtS+9mYWJh5mVWruNPLhfN6tTN4M7Rl3P85AvXiY6fqr2+RKuZwgG5KNJyN7TzuXsFwjuc2kv45Uu0uJPOGHGjMuwy0E/Fc+wJ2D3Qtjp3pepp/FFFlRmYCd47FxjM2Z8pRieew6HW1/61Xp92HdEJMIszPCcUy1V1YhyThyCaDNXdWYCoKpJhJk9FuGJ3Q1Ak/PwLjYGK5wiFg4+HUSR0LYEtLubmzORAyln06o1Srl9xhqgwEmn73x0dHOxvHN9uazrVE5RVrnJzaJp2iblJqUkLE3T5twwc6QdfKuHGNGN1brpuvV6nVJS1a7railmxiCtvWm/WLTtIjdNXm0KH9y4+f0fFGdUbVWMjv75P/1H/+xfzKEIZ8yYMeMFxkxAz5gxY8YLiW51/Iv/8K+vLxbXD5e0OYZprcWZ3LwUraruzkwwV7NaOtPqrlY616rGKaXUNDnnQThDJLlp2kVKmUWIxB1gpoNDliSAm5tarQaWh8cnf/HzX7zz/kfVEPbRg9lfSFmCznC88sqr/+Uf/RExf/rgwUd377bNtZQXFk6Gbgq4w3QgW82MeZhr9aV43wNQ1VoraLAzDPZZ1YjAzDE7iliFqhrstKoBHt6ItdbNZnNyfLxZr90MA4f+1WEvEfxF4OFi4k8UJF40zdj98wmS7pldmvEV4am9/WJ/9qcZsF9x+FxGZH8VQ/0JlPcLjWdYDJgxY8azYRhuRGRqfd9prU3bHiyXwly1ugU/TO5OzCIyvd4QCRHlnN1d1cI7GYCqg5w5/C5gY5SLieQNeXISAVGw04NgGhHROeIFIuWkVWolDAbUFOGkHTCgAivHUdGjjV47PFg07GtvFm1qBBSvX2ZqpRQAKWUREZHICD0RTw98T0mIkHNu29bNzUxLcasEa5pMTGaWEnu100ePvD2wTaW0YCwA/drba8aMGTNmPE/MBPSMGTNmvHh459/8y5P77xGnxWLRChXd1H5Vay/Ept73pdZq5sJiaqpqqA6DO4k0KRNzSo3kzCyxbdKAlJvF4WEIZOAOd4Csadzda2F4de1LWfX2yb0Hf/XXv3z/w7tVd+XEW8YniRweLN944/Uf//hH77///sd3P/3s4dHNm3lJuSrUzd1hRiA41BTuqhrWz4BXVVUNWbSqTuwzAI/zgSmku1aNQD2D6sccAMgBL6WsTlePHj7qNhsM8ufhu68Q06xuInSc9p0w/rUvi71f+pn/XMzKR9XSOfhXTTD5ngodKW/aPYN2iEoHELNluG9vZF9eIAwU57m9yLST8/aiF/+8Cp5GoZ5r1r3lPJPPs3kiPwN2LrdlFHaK4Lhwd5fXDxGNmrXdY37p/X51uMoSzjfFnH73DCv2btF4jo1+9ayeWrGz4/aM7wQc5lqL913XNM3h4SERrdfrTbcxw2jl7ABVVa1mZmwerG6EHJwiMIe1BRwsAiLVCoCYmdnUaqmShEDO4yYyMyImEcDdrFYlAoNYGMzE4gbAopAYl8QV6IDjoo835XduX7/WtMiU28wCs5okiSQgYkRrSiRCInCnWGp0D3GAiLBIcoewtO3C3VW19j3cmEBM7lZVU6ZqVMqGUtskXpuSFEn5X771P/5Pb/0v31yzzZgxY8aML4WZgJ4xY8aMFw99zsvSnTbCBPTH5fSzfn1spTAYjloNIBh1RUHMSdrlosLWXXf9xq3F8hqnxkAOzjklSSLiACWRRUNw1ILNGnC3Wh8da9+plcRUSj062dxf8a9+9eEv/+ZXn9x7oAaHbvmAQVTjy2X74x+/+eMfvXnnzu3/8Bc/e//Dj7vixSkTK7sq1Kz0VZhykm5dtVZVbZompYQxQs4Y4V2YyeG12uC5AbchGDwBZBYBc8BE6jBzJjK1mLHVvj89Oi59F1Hdg934wpbJdGXOmvaxJ2NQRAz83pZjoYtsy6Xs5Xni2ben0c7/z197IKbj/09laM/5Pl7AaEd5NoldIrsmxkASGwCKP4PMdANAnAhuqiHscneHjS21vVfi0ePFbYfaJiJyGHyqYRqYQaKRIL6s3fzsrU5JHOA9CYmIOYhZIsa4vxkgMMF9KMMwzzYAIL5AUk+Mqu38eaEk29P48sLvnrlt1NjK4G4YK3yslZ2CDTe7W57pszExiFw1th3AnOLeTR0O4hgJOxYxZ6nubTVi5/i5a+3eCC7XQT+V5N3LmV7253PHF2JUp974QtDWdGEp47ngKlk9WRQ/nfPlA8nOmPGNwt2sAjDy05OT5WJ546WXTHW9Xq9OV5xSzo2q1t76WhE/feYAmDnlFG84xBQaglqrVu3dctOwSC0VBGLSUswc5lrUq2nl+J0tpQqz5YTYZ1YKMTGTKBuIJWsYeMCG0ehbEfRJVx6d9tIubt5sW1sQxzfWtm3btiw8/AiQw82hg9+07LizxY9IXCnnWmot8JTji77vnNAulim3TtKraVos0Zw+2ij84OZh3/ffRIPNmDFjxozng5mAnjFjxowXD8Z0eniIUrTW1eZRtzl1LRR2GE7iIGcwC6eUclos0uHCCMta2sMbuVmSsVGcIOE6XGvVvvR9b6XXbl1Xx7Dqrq7VVE2rlb6Y9ZY//vj43Xc/ePz4pNYqHPRz0F4D8UTui6b98Q9/eO3w8O7dex9/cne16b/36mu5XZAkdlASMRdVmDHQtkJti1FUGqIeIpg5M6eUzFTVmLXJWUS6vnd3Is45AZCqIBKR3DTZYdkJUK19R6uu6zZdxDZ85qqmM5wybY/sMr40eiaeZZRpPMe3HDHRdHwQBhF2k+2KheM/k4/jDq/HmJy3t+XcXvpsufZ+AYQUfIf93G7K3XKnROdYqOBeg5YkczfV4GWHxQeHuTETMw+qLIcIAVDVuJyaMnManCiJmEa7yoHYFWZzUzVhJkIEoqRISEzEka3DQwhvg8hqexdjbfkZipaIic206uQ8Hkw2QOzucBszP0+yx80RYepLw73xMJ0mYiImBP8LikBPjjPdZ6pLdw9WmKLG3H1w4TQzplhZ2aM6jgWZqQBm5j4t1QzDUFUBEJOwmHnshABgUTDQ5M45lGjqEURDeUyHMJ5mE63svu0YPKrAB39POvPB3bd68bM3vsNYb8fFuDQyDZczBdtRx2N3JI0HRy7+zJpNdMMI0XWuMb9m/ez5p8eLgqvoz785fLtLN2PGleAA3Gy9Wq9Xq1qVRdq2XS6XICIWd4hww427E8Dg4YEGsLBIQyOE2bLZuF2sbRuMy4QsSCIAti8f7sKM0b+DiYTFoUA4m5GLQ8n97DN1/N/Jqr/74PGDh0c30uENqXAlsmEd1n2xWEialNm8fc/hcYGUeTjkIBqMQbz1JAw31bLZQA2cGpbkJOIwyU06uKP0eN2fnJxma//kj//4n/zpn37dzTVjxowZM54HZgJ6xowZM14w/OIXP7WNQ61ps5f1anXkWoVEchJJBOYKciKwsOR2kZcLWmQIuzukAcT7GhFp4OpVa62ldKXvS19q19XNql8fmRWQkwgRkflmfWokadHevXf/nfc+OF0XczDDDB70nA4MFTMfHhz83u++mVN+++137t37tFR96fuvdH0tajGPIkdKoqXWviyaNqfMSbquq7WKSEqJWVQrMzc5d31vVpkhkkWEqTqBWYgF7kROzCyJSEAQcgLcDER91282m/BPfLaqngjZ8cMwi9rlasdI8jR+2KYdiWaaDkStD4eImOMzgQbh7Za13OG5x3hC7iMXysTB2k1uC7RT2jHd8K9dbnr7MWaAOyUeixe2GORw2pZhYnMd7kQ8UsxWq8aZIgIEAVpFRCSpVjMHKOUE977viBlEtdYk0uRcao1vVdVtuEcQckpqWkrJKYOgtYokZqqqwiKS1AYkEYDMwrBldBIXVrWh0WkSTYeOWWqtfSk5Z2GJW6TJYdwHRvsiZxk8LxNUw/hcfBDiD1Nsj24oolVBFLfg5sRjLW4dYOJStr2umZmxCNxVjZndobpHWM5ESSTk2GMdODOIiYncXE3PENBqqp6bTESqIYsmER7uKvqnY1JME2BuahbWPDZW48Tixi1LON4MO8RBgJmPBL0HXRKJxq4z3vxo5kFEDoLTyCpv12R2NgxM3XKnAhkAje2zI7WmaUHG3Q1upfSxtWKn+FNn3itGvkyhfPH4BX79Urwoqudz+AYsV2bM+C2Eu/fdZr1erVanIGradrFcmrm5q6pIypLMjIEkKaJixAJqEhljDQZxDFVVVQeapsH4s0IEZtl73XHVkIioanVXJq4gMx+444upgNW6v/+53/3s4Y2stBTTnlxzYtl0OafDg5KbnJIQgwhMFL+AsZGGmYQH0LiOzQJmbheNm9a+JyY1gLMTgZiIXBrPzevNgX726HhTaXVg7forbpYZM2bMmPFVYSagZ8yYMeMFgxfDgtOaX759U7vjfo3ULpOklFuQiOQkOTgdlsQiJERWYAaRcnqqm95KjcAvgFbtS9+V0ps6uZSwG0Q1mAJuLjnntkn5QNKiPbx9/+HPf/32u6frXo2c4XAYnIc9l2S4dn35vZfvvPbKq6Uvv/7Vr4+PTkqp63XXl1qqmoOCI3YvXd9tuq4pbW6aptlsulJ6Ik4pSZJaCkAppVpKrVVNc96wcN/15h5xCN28VpUkKaWcW62qWsnd3Gqtx8fH3aYL6nCcTdHVmJXzJxMxCxMEId8ZVNqgC8D2OGKWNbLNEyENwjQrAw+feBKfxvUZPCUZaGmHAxyqIeJBhrrz7VjULfccdBvRJD8aTxkTxilDAUYy2sf0uwmDFiQQx5oEkZv5SBkyk4gQOBS4xMTMo/yaQHDzUkvOjSTRWolJRCY5takRICmZq8NzSqpaSg2Ru9bKwboO3DcH+WlmIkIgNY05dt93Oee2abq+N9ULThogonDPjIQAiGTQIRPFf5mI5cyM3d1qrXADIaXEIgQ4wcxKKdGWpZQkqWnaru+ZaLlc9qWoVmYJX/W+9AQSEbXqbpNaeCRYg64lZja3UC5fNAKJVBxUt4iZmllKQkSA16puRkxBUhDg5g5ftEtmUQsFNGLLtpklSdGuVYubEUE4LEQ11hrMPSiCWouZMUeoqclH1HgQyLtVDTl2FB3BRJsG3zttj9i9GTgNVvODgHlLNU9LJxhlc9EMYZEyLqLsssBbBXwEw3KrJyfH69Wq74up2o5pw7COs5t26h/jKdiPp56wFy8Wl+vTahOAF5M9nzHjhQKh67vPP//s+vXrAFSr+7irLPjl8U0g1v/SsEjPsbgeB+NHOezUtNaR82V3U63xIxU8dSQ59ycTgSRsm2J52Z2mJ2VshIpAhRXozB+erI/Wi1sHN45Pj6zvlouGAMCYH7Vt0y6WRPHbQUQkzJJSSpKyNLlJOSeJH1JmdsAZEAO5gJvUcGZOTTNZeBmEcnP72p1COPnkQb35kPvmG2qqGTNmzJjxZTET0DNmzJjxokHhRXOzPFgsq63S8jBJcM0JziBmTnAnD6aplHWn3cZdnci6aqVYqaYGM5CZlap9qZUgWZaJOAARi3EAACAASURBVC8WaXGIxEZQYsltygtCMk/V0uePN/c+fVSK+rAHHz7pGAECbt648eor379+7fq9Tz998OAzELXtQiS1nFL2qhr6RLgLUU6JibPkpmmYuWp2d2EJa0NzJyA3WZKoWWzsbFqalDtmBuKcE7MMDg7mEZDdTfu+6/tuMgQguiL7HLigefQdz4aJlR3ZY6at1Gd7+CxPPamdaUo0JRzNNtwECJU4Bwc9ip+3ZPGUDJEG09cYPR8mMjmY0i0FvqN59snQOYozsng+2hyMiUZdatQDMw+MLUvooKdKARE58aBsGqsp5JTsOTcSM86w5BjrwQFJw+ZcHm+ViMMlgwiU87ibWOAxCSciDiWvA8zBwEIkEbHF3l7BOe4vKopFcs5mU50RMDCtRBQd6LwbBDgl8ejmg1d1WGeAWOJUSYmixxKBaNB+ExOzE6n7VCAHiDmlVEp1V5Gh647S86CIfaRZtxgE18w0/Q/OhOhn7u6oBiRmlpRHpj5uGWGk7YOnczDsE9FIHIYkTiwg0NgD2EM2HvnbmKEN/wwUhbvDRGMhxG2kqN3dbSSox4qmnV4RCzw7FiDYLp/QlmXeteAYVmBi8/i0uDOkjAY2M7dqWkotsXTlbqS062DzrKTwCypnfgZMQ+O355ZnzPim4H3fHR09zjktFsuD5UFVrWqIzSHuLBKvAimliT4movFPnezLIrvphMh8Z5lz+Hv4vRjfo4Knjud2sNgp5wq1WrdFHB8HBnRq9x6evHx98epLdyAtZzCLhAGVq3nstgmbKQKBiSSZMLEQcxfrpylxSpJyjl+lnNc0vupITm3V2J3jZiQ5LcCLkiW5Vaama0/feusfvPXWv/0a22jGjBkzZjwfzAT0jBkzZrxI8J/+9L1TO2m4TU2CNU12vkEcXCTM3NS0FLjHDGN9enJ6ctz3XS29a825ZZBWdTM4RBxkRgYilqZpDznnZtke3jjgNkFYHSSZpSVqT1blk3sPP3+8efhoHe4Ag0fArmeu4/bt26+99lpumr4vq9W6bQ8kt027lNyAqPS9ajVTmAlzklRKYaa2aYOLDAOB8FWIDaciQkSqvtUujrSTmdVac84A9V1fa3I3Bkrp11ar1jB5mGhW/yIM9BaTDNkdNNkNj0bDwXxNPhuTZpPIJ1o2vuCJfhtIvcHwGgQMBBmJEDBwzAMNOFHF7thRVe9wbwgqeltgx5ZFHSlgP1MJoxnxQGITbJjvTdzTwEJu7Q4mDjpqYryDgeWcTJe3WtazFOqgn92y5TSSohBhIoSca9cxw91DW92X4mZN09ToEpyCdA7BeKwMjNPs4cNIcmI4AjhQSsk5LxfLru+0atSowVWNmFnYVIkoSRobeGhUYXKCu2utFvWlRkDK2cwcnnN2R602XFgtZODCom5ulnMGUGt1uAi3bRMG5U3ThmycmdwHD+iR8qep8ABKre4uIsHjAzBTd5OUCDC3ruvdPacUDZObDIeaua1NTc0G/5YhrY/uNJRSitqOFovC/P/svcuPJFmW3nce914zj4iMrOqu7pqe7pmmRtALAqi/hksB1IYCpK20r720EiAB4oYEuBvutZLQWugBiJAIjIihONNN9nTX+5GVmRHhbnbveWhx7jX3yKohu7qri5VT9gGVFeHhbm6Pa+Zuv/ud73AMxe2o98PYKTOCA6Jb586wEZDRsBP7cfHzTEYf8BS2t4vFDT/yyAvdJnJg+J630TicfEQXsypjUWHNdpWmgjllZkZCUHzMnL/qReByGF+apl8va/NvqMs9dYnsd+3a9fuStHYvcn11NU/z06e3x9N6WhZiVjVRo0hYUo8uza21eFXOGUchjo85TgBgZh/RHDER7tvk3Pg4jy9XABAgW1XUzM0QiJkhZ3CpUh/VQ+AZQH/w7P6t2+t/z2m+flLgUEBLSTlx1JoggLn2y3F8rLiLqjW1iBcBZ8acU5kmt4vPbnAETCVP0wwOrm6i5TBPN3USroKg5mDPb55fy5Nv8gDt2rVr166vSzuA3rVr167XSZ/cwk8/ol/8VK7njLaimzvoWrU1bdVU2lpPx1PExKpZq02kMVFxMGQCJC5cEhIhEzI5uqPnPOXpappvqEyUiFHcddgz0aoY0Afvfvi//u//16/efU8dzMEx+uBt0A/cwQDe/uHbP/nxTz759NnHnz4T8asn11QmdVC1MIRmzAQJPSICoSQeeNUQccrZI98WMHG+OszD2OhBopvI8Pl2GIbEgHg4HFTV1MD9+efPXt69rLVGR7ggrtbbun0RpnzJI1/wPw+o6lsDOQhbdCzdgu4ROEa67QWIBoiNBer5AcMevOVyYC81daBz8MD2p0eRxMMiut0UPqZgvqURYNwuRpe2jY6fbVAXqR2XoLu7ojYT9HlHIMCjXYVIFz8jEsa9JV6wdXcf1nW6sGvHXoBxP4zMtLUZjE6DRMREogoAxL3WOAgsABgCgESSBhEReWRKMHEQfRve2sTs4K01ZiJiVxdvJ7PWmqnFegcrl9a8eoR+tFbRwc1FBbsNu1uke8Iykrs5eBVVUwAgA1FdlzbPEyK22mJdamwvQbQaFGnMhEqrqIiY6tI0RkNUQWOUYENPw3D3VoWIck6ucUsPqmaxJugIILXGsNTIwiYyBwcFtYDFAKhqrbXYXTpOho3dNhUMpxohgJuqI3rvEnkeGYQwmvqNWA0fVug+kYL9AMdWwxa+0ediYHjqe/3EMNieyfM2Fvugoj62xnM6xiYeSdFnb1/kf7i71LYup/v7u3VdVNQDeHSQ8ptA1S/90yV0/qoRHK8TwP0ibt+1a9fXry3mphe/wMPDMU/zzdM3/Lgsy4qEZq5muog7uBj27n7hLMZaa9SKBVyutV1M7Dm4h3MaES1QsFl89RjlYgYAaqZm8U2JkM3cXImIOXFK1kvWBhtGcAB1uBf4fNVnp+UnT+fbwzxBKzmlzKM/rfcJxagDAzdXB+tLAcQoXwPkxKZRycattdqaiEpTgOpq2kya8Cp8Mn4hK89eVbL/cPnDE+4x0Lt27dr1WmoH0Lt27dr1OmlJ+uc/4Rv04tLu78DEzWRdpS5SV1CRWtuyCCACijsAEmJmJmYHolw4zzzNmDMmBsLgR6XMaZq5TJAygLdI6lABB3B0o9Ny+uUvf/V//J//5P0PPo5w2i0SAgLHOhBhTvy9N58+vX363gcffvLJs9Pa0kEZpYqqr+5ABAmBEQjRzcw0peQOTdqoxMzmZqpmTswpp1EbCgGgRRX8UUCBg8SNTjggpcnxeLx7eddavUS3m3/6sfDiwcdxAK886/LJsaxx3+gj2Bp7Zzm4wMDdV4zog0dv7PkccBEozh16c8gzi/vi6uDmCsUv+fPljumbhNsCxyae2fPFLvFBDnFQwrFEgM3X2rc6zNSb7zhyREDVfMwT4HBduXtkSkLERg+rLCI2aeYGgIkTE7q7qJgpc2JmIlRVM+8G8osVIJQw8KaUhkFefQDoQNsAjojWLWNViYgoeuXVdWPfMRlAgCQqqmqaCSn8tmZWW6POP73vh24TxnCiRxQyOLiam6toBQeAVhszI5GpRaKMjuB15sjPoPA7R7NNZrax52NwGSpERE5riKgtxXEzEE4MgK21mOvQ0QfSzYl6g8LY7d67GrKZa7RHRASiaGDpI2FjGMkRwxytEmNTR7qoqQIYIQ2fcQfKGu0gPeYYNsh7nmnosz99wIwh18n1eS5ihNC8en7hcEzH8oNc4whr2U6TWLJprIu3tS6n07qurbZxoH9HlIoXP3xV+vz66W+wwXvXrm+j3AFgXdd1WUyVmXNKp+UkIrZFGsXlG3sRFACaGyEyUSBmETnPSztA/+Ttn1Nu7r2HBNoXv+M4IAJzMlMz5dFxAdF6+VCQb3ADEICTwotFPn55/9ZNdiSVquzJkRLH+iBFWFT/8AewaI2NQDHpaxpTsxS9QZBYRFsTMQVAItImypZzAWAHtFYR8kz5iKDNi+8x0Lt27dr1WmoH0Lt27dr1Oun5pGgtpwL14f7Zh8HvpIm2aq2hGyHknFXV3Ik4lamUKTNHSHSeDjzNPB9gmiElUDGpKoLEjtDaCm1Vbe10r61aq22pRIl5/ujZw1/85S/+yf/9Zx9/fnKAqMAf5fUdiCbmpzfTzfWBmD/55NNPP312d3+sRpSKOSx1VVEmyoSJgBhFWl3rVAoC1lZ9AOho5s7ESAhM7g7WS/BpdM55RQ4A2JNtl+PDs88+u7+7C1PPV9GXgpcwalO0AoJB1Lb/u3cIHzkc2DM6OneLF2DgS3TcMgNGaHT3OAfXM6fNVowwOC/C9uBAeuY2MDFsluhuJiV4xMu2zGnsN6JbigCe36hj9HBFDdrXgfUFuI7VwaCH2zIBw2buw2oaLnCvrSFEbCUgEicOQBjEmZi6DRkAsgtCizkP8FyKSA/AMDNVyzkTkwwHNCEHvQ1L7/CKo4J43Gy7IQIziwgiRhfBbYFmFqNIVZkiNtoDPy/LwsQlpaDYrTbs5uxurx35FZZzZiLTDgdOx2M0IVyOJ1VVtYDj7p5yAobT6RR0Xk2IcColpkxarYjIzLVWc2eiUgoxq0Q/P4tOg+4wTYWIVK1MhYjaWsNTFhXZKaXID3Ht6xRcXkUQEzMx07JWM88lp8REUGtDxJQT2JkGO4Kqdi+2WyfR0tydExEROIT3nJlVRFQjsuOSzXpYpe0i7GUbb9FAcvDn8+jcQp834z4AbPi5M2g0204/vxjb4O6mqqKmJq21talpZFWP8Bno5+Jv6mJ+nWzLX6PiVHq1A+auXbt+P9qmyc201vV4fz/NhzeePn354vnpdOqVQ4AAHDFeANBn+9zALPpLj6cNmYM7Mve0LhF3A0498Ij51eubOyAQiZu6abQIjgbGSP1a2+umHNShArxc6/ufvvjRk3IFye6fHebp6vpwOMzTVHLOjNS/D4EDYsmZOfoW0DZ1HunQtVVRBSCORibju0dbV1dPaZJmtYkYCJWi/uHDutTVU/5v/qv/9L/+b//RN3KIdu3atWvX16YdQO/atWvXa6N/9rM/VV0N3A3qw0tdTwAAxGAOyJARiZAYOVJgOZe5zHOeSyRDIBJS6o4UE1+b18Vada3mLmpV2rourVU3qetS1+oGZb6Z5tvnL15+9vz+5b0s4gpRSzliHKLQ0v36MP34R394++RGW/vkk09f3t8DcWsKWh3JFcDBRKtrBQMIOuzH0wJn466L1iBuRBo0N0jW8GKOjvCv+H7DF0sIDrWuG238rYSXODceChOlmY1kXgdA8M2c637ehLGUbuwM87B1AB0pJFv6xniLnmjAryLwSzbXnaXDQBr8elvHYaU+r3a3PdP5LxAkP3hgX4luhe3hGw4APgJ2z9kdsK2Vb8fdI1gjfLJR4EuYEHA04gNmivcJDyoREjE4mbuZqHpOTDnHzbQDpHlyyw7ORA7gbhF5GS4wcM+JwyQ7ug7igOd9cqCj+dEHEQmbNnBPiR3cINY5MH3wSAQEJMjEnMidEcnNRFspJXFiJu+7C6zHg2DA3Sa1uoP7NM1TLmslQqJE5ISMpVt0Macc4Rhlyt5bKiUiRO6OMmQ0MxNLJTm4NFmlsqWUUtjqmVMmYubY8ZQiHtw5kxmYWZkKMTGztBb51EhIvV1kP0kd3RHylGEEngD4lqdsADC6JgIAgMXwZegB35zSGAKxx7pZGQmjX+b5tOjni41zaYuzHtbm4YwGAAC6eMZ4fszbjGmSi5MgGnE9io4ZOMbdXcUQVaBCizxTH0P6MZr5yi7mS33VF75+FPtiC7+sxGLXrl2/H5laXevd3f0tMXEq09zM1DSnhBDlO1u9EgACE5lqqy2XTERRsDKe4O49DssBMCV3M+9fn744Mx9fsIgp/oRE4ObRJeHychxXdgQAuFvq+x8//+M35isv/vDwcFzLwzJNOZdccsoll5JTSoSABIyYc845p0DMACXnlHJiAEyJmThF5VPkMwHAlA7xYaOqs7K7K083PC2fvPjsfr3nwlh/f8di165du3b9nrQD6F27du16beSkbFPzB3Bv6xGi8p0JCRnJiYkTckbOyIlTLtOcpkyJ3RpEGrKBmEFbrTWtVZajS3Nr5tpaW2td10VVUuJWW2vCKSM4Ej+/u//s+f2xebMLeAwAAOiABIhwc3397/7Jv3NzfX18eHjx4mVrMs+HKm4OGI3diNxGF5pw2nKqKgAQndPAXcyiRR9QZ1qI6Bj50gAOYrplBWyKMGYQMLO1rnLRvf231avwZTQcxOEZhgv8C2ekjBtSw5FdG8Znh0cd1C4ClofVeSuf3dYh4pQHu9vYGwKMOOmxshce0u3VOPKmt+SNTroRI0ICg+iNrAyIe026eM1IkobNYLWtBjMjEiCaqpq6O9NIwwh3EzFchC3gcK+ramtNVUrOgZgj4jnnHHMNHQ6DJ06xwBYRz0yIhBB2WGYmVX3FmLyFfriDujmYuyEhAjFCPM7MHf4SMfUY6R5abRZ9DkvOxOTWHbeUyNxUBdzNjMxabW4a6cxlKuG+R0SkEoc+ci3C0S8iOZfYUjNDhJwTRg4mQsyX5Kn02BBzJODE5OTJATDnVEqptVcJhAk9YTJTc8qp28A5UWRiRII2M1NSrBSLJepP65Ex7ilnImImNHQnNAgD/oUpGd37AhHATGPAsTMSxNjky3mKc9ByjxMhpEdG/S1lPMzNSGMCZgzZixyOi0XGArGfcwiPWxv2OBEVE5GKJKIAi4/pki+bi/rtGPR3xBR8uXN2+rxr1zckd2ut3d/fH66urqbpcHVlCFVayRmBVGw8LT5PIacsooDUi2MuAPT2OXiu+HA305g2NnsVQZsqADCzsplyYnITdd9SsxwdI0kfwRAc4Fjl4+f6/H5960DZSFSXtqS15pxKTvNcSim5ZHAHNzcrZSqlxCe+ux/meSol5QwAiJiSM9kI6wJETykTo4MnwpSIGJ1Z0vT9dvVyXSd88Dr/j3/v7/3nf//v//6PzK5du3bt+tq0A+hdu3btej30p3/6p8dmh6nNaUIiByjznHPhXByROFPOQBk5AWVMDMjopiLr6dh0jVACb+oiWtfT8WF5eGjrQmCJwd3FtIlMpczTNM3z7W2ilDmVfPUGpCfP/+nPP/r8846xATpfAgQwQDBzdHhye/u3/5O/zZw++uRjUT0crq5vn94fT6JGnCIJ0MHcFEzBLWr0c1FATJzClKqqwa2059J2t6aIRjP3dV0AkJkvd467u5qIruu6rEttbRSp/i7abJk0mByd2TeeTcQQRt+O287BANHUrTPogaQjlrHD4x5OsL3VWOdRZtsTHDfAd37DcyErQM/RjWWeETV0Bj1MoBd/GCsDgD0h9+KvBNgzQ7bgBD//M9j7loWCnvwRQuz99qyHRFv8FYn7zbCZTaWoWcQ3w4iETimripmmnJiZiVqL5Ic0z/PjA0PhlhKRoLeX99VEmFJS1WU93T65RoDj6cTMKSUfCc7aPfKYcyGk1uo0TVOZ7h8eJoBpmtRURVtrGP2YModRu7Vqag6ukwLiVEpQ7+vrSdWayNX1DA7Lss7zxMyqljPECCWinPl4PLr74XAgJnBY1zWsaioCiFeHq9jL566brTFzznls4PlxB0PEaEIlItdX12Z2PB5jY3PJptZS27zqkVsiIpHOOU0TjmCW7mxDBodA5DjaSLpbT5Vx7R5oopi2iAG/AY4RwQLn4b+NzNBjb38H0BfdCGEbmD12fHQ5dItLDzH22O5t4I8Fm5mIppxV9fTwgOf4jVffG76aviPcuWtcgL5bW71r17dAqKqn08nc53m6fXqbclrWBYnAEXKfTHOz+CAmpJTSNBUAQIR8OV8+rs845g63wCOAL5RrjTlgZo7MK2YyFSFaVOLtohztvHzE5nAvcFL0dLi9vjFdTVcEm0qap6mUlBITooiKNGnSmq5rA0CR1lo7zHOZckopkpqIOdpaH+Y55USEpaRcSp6m+DaQAM1qM5pzKUz3DQ/Hm5bWb+Co7Nq1a9eur1E7gN61a9eu10NvHeyvntF//BP/wdtvUV2Qn06ZUiKingyIiGCgra3rQ3Q/d9FW11pXAzUwMzU1VzU1U2UCnAsgEGIgwAQ4z4dpmkopRIycy3ztNN8v/otff/gvf/WBjATWRwZCB0R4440nb//oB2//6O333//g088+neapIJecruZJ1AIxE6KDgTshMJGILOua3IgopRyAT9WYmZlE+ruFV3SYmn0qHPZXVe09zADcXNVPp9O6Lq1Wae2CPPlXREgRLjCCLeIhDL9mB2oX4bPdBY14Tta48EJ3Jkyb+fni8eH0fBQ+MGgdjrZ/eL5rDDK3Wafdt3DbvlawhWqMxeIFf9uI8pb7cU5CQKQN/0UaND561XmJtG3vec0JEWhj04BAHhW9gIicuXNhJDcDN0bklNPZNk7mBg7MRJTdaLPREpCjEzGMkOzxju6m6haoNBornXNHCBGBCNOIiD5MU6xMn/QA31JQomshIbqqtErgRMSEKo7gcylNxVQgxTYCI0cUcsMGiPM0m6mImGp/I3d3Lzkxdf97rMW6LgiYmOdpCp9yGMajZRMxKxECxMzKMAojAGBOAOhmTMjEY8DBVEqQ6sjl5BIOZzrMc7c7IxEjEwFEUQGZmarS+QiOoBj0MUgZHM0NNiKMcb4CADhw98VTdCPsA6+nfLhbd833rPZh3n/EOi4DN2Ie61wKcD7Ztghyd3I08zgjRvDMNvw2moKAQJQSg3vOhTmZbaUa2/j9StcBf2XNvztyePWYfB36ju7MXa+bfsOB+rvP0HzJG7m5tLaeTsuyZOZ5miDoMAAxx2QnDhNxLAMBAx/T+H7hvSOrxnsgIhG79wKhuIa6u5lt32KiXUGsQ68JwoRgrSVzja62j2b0HcxBwD97+fDyeP3TH/0R6WLtmMgzY06Uc3z4gpWkkltTREJiIlLhypgzI4BUiU0wA1Ux1VplfBuJor4cn++JCXKBfJB8A+qufDrckTDs2rVr167XSjuA3rVr167XQ4X1P/qezXN5883beoeerUwZwMAMiNzMRbzV9eH+7vnzzJiQXFSkNmnIqGCi2uspHfM0zVdXnLIhmgPlTKkglzzNKWdGNjMHSjdvLKt//uzZz3/5/i9/fQGge1Vm/AJI+MO3v//jH7999eTquByfPX82HYp7AveSM7OZWU5ERGaIhIkw57LWtamQExHlksEtmrBF97bEpKpqXnIKdgtuAD6VzhVra24+ch5A1Vpd3VRq094O3n9j+oxf8tuZcY3cDCLYaO8FgB72Z3gEoAdq65G5W/LG4HrnXMVuMsYtYiAw8LjHxAg5jsSD2PcGl26kHoSMuP0I5/iBLUljGKW3F4w72M2hOqj0yC04m8gfG6YQcBDSaE504Y0aIb/u4G4RBRE/A3ike0cHQiIauRwcmSyImJCAqNZmZjHICImAotNdPAcRwN1UzHqsBxKPdY+cFlR1dyBmUwPEnLKZ9rwO62bkAL8eHQvBVZpKQyQEl/gZIE+5SZXWBlEFcKce5N27PUbeRa01p1RyPh6P7pZzAVdVN7dA0W6q7qY5cSKwZV0JkJndHAnQnXtcd7SDAiIKYMBEZqbSevAIUSy3J5YYqCkiMidXB4SpTAHrXS2maswUARKTuAMhJg5HcQAIZog08202hRBHfUIfSLFjkcakhVmUQFhEhHacsTERBCSITPZHaRp9LI2R5ps7/mxjjr9YMO5wgts5xQXALDzsdp6/iB2GDoAEwJxTKiklFTGER9Dkt0ze+KK21X1d9OrV4iu+5GtZgR1A73pd9G8cq1/jZWRbGo4iI3s4PpSX0+3tbRkJTu5AaSvx6Wn4Zr1JbFwkYZuNHhPHWz5VfK8IH3R84JupiPZPwdEaQVXPK4eYUk65mJlKBXvc1HnUQ336/P6Tl0/46smME7U0JU9ohJ6YmJCjlQCgiJuDQxQnSWsrEZtZXRszE5I5rABqXkXdXE1rraYKiN0iTYRl4umarqtO1yBuoLXIO+/8nXfe+cdfx+HYtWvXrl3fhHYAvWvXrl2vh25KVcKUrgGcQKW10+mhtVWlMSGYmai2KsuyHI8lcWZOSEQwTcXcmHKZCBAdwAzSVPI85WkGIAXP04FyAS6UCxKju1YxQyxXy/H42ed3z16c7k9NDNAfm+MirY/op3/8kz/88Y9e3r28e3hYajVzd3WIjnNmqpU5QFXU5jOvTdqyrGFr5CajDzs10SB87m6qp0V7sIMpgJec1cxURRUBU8oAoGq1yvF0Oi1LN9/+ptz5ryEjl5u4kd0LU+SXE+u49/OA1mcnNHTjZo9+hoEZ3belIgbJAwSAoKSA5+wPiMZwI+LAwQk8joUjeBBg3Crnh5nJNwt1sDeHPoOw2ZXjaPpluiT29RvdhjZAfcbbjwFcB6c9THp7fvTcU9FITzDvqD6SJfsT3MyEEyOAiEA3efeMElWNfHMAdQdwYiZiai3SkCOeBc2dHAHQzZlTzqnW5u5EHK0Dm0tU8UpbmVOZyrqsZl5KWteqqjkxUUKKDGhzNUR0h+NpAaSUSq2ViVNKImKmZp6ngkQv7u77DASRmh2PDyJiZrXWLVd60QXAAyK01ogYAd291gYgIi1GRhNBwJyTmpn5djqklES01hqtmrpH3fzoJ8Ce2hzEmZjjV1VxgKlMiGZuIhUAc84RtTF4bnBnFBJ3x4vRAxezH96H4hbh7X1SA/s0iY+5lHg6IRGRupgFqMdHl4tx9YhFuF8OJI9JlBh/ZH1WxUYGR4xwHzMcMKoOumXffTNWM/E0TSqiKg6vpJ3ixQ/++JEvXjFeI8T8r5e/es7u2rXr26JXv4E8PDwg0ZMnT6J+5XRaRGQqMyK62/EoKaWUWNUiZig+Mc3ikwNy7xm7XS23OcL42PVaa1zP48EtEvoCT1t0EShlMjNpLb6d9C8f8ckAYADPfcZjYwAAIABJREFUHuTdZ6dfffzsrSu8YXHRqdBUMjIxY0JKKROyOSAy9CYQYlJyLggQn3rxIS4qTTUa2rpD1BVt+U5m1swbkGgT0XVtuaTjU8p1Rxm7du3a9Tppv2rv2rVr12ugn/3sH4g2VkW5evHhe7gcvS6urdZVWiUicDdVUzUVADdwRaBEnBIyMxJx5lyI2QnNgRJz4sQc0X4RKwAIWtfWpC7relqbQHnQv3rv43/6//zZx58+q2KA4JtPZ6DOlOjqqvzoD95+evv0vfc/+OSzz+6PC4CZoSpEukK3rZ43CDEyW63fYFA0NMfgzgDgOSXAnk7roxEOEdbUTK215mZIlHPpNydNHo7HZVnUX22w8xWFA2V1jDwe74hrMOMLR6fbMIUDADgCOlBQYuh9exzAccRSbM8cPGh7LSGCgw08TNAhW1+zDm3BwGjDx2Mdh8F5kMMBEYOK90CI8d7brSai9RAEH92NABAizhcQYASPwAhaGOuyHc8B2aNQFzt3RItFoQwe7W4O7lsSiWnn7CwMAK22QK60MXczAKwteus5AIgiErTaEIFTjrZLvS9lly5rVRV3oMiWMFdVTkxErbaU3BGrSMyQLMuiIillZkIid1dVUU3MkXQcR8dUEZVaE5E4OqspIppa3wE0TNgOaiqizMTMxOxmqrY1e6QRYYyjfZ6P3okxEyMRx0lERICIa4tAaqzIPXzGwkvOKaWUgiCYai6FCEVUVBBQHQBQRGpbCXGe5zEZZJ3wj5EAfYqENyddePrDJe1mRBDZ5dtf+8jvo2AMfnfDYPdxzo8OhDAyZPrQwW6TH6eYI+DIlXcAB8fRn7Dj54gI6bMx2Bl4P6/6RiCeITkTjwD2XV2XoP3rsoLv2rXra5fUui4nEUk5I5K0tq5VxSn6EIhEkZiJxMcGRZISkUpzM0kZL+u/3BEpZntj+T5s1GYG7jAaHQ8hgjMRM6na+UrhfnkNCQD9IP7x3enn737Qvnd464qL1ynzNJUpc0kpM5XiiRM6EkNKmEtOKXnKOSfevhY6Olh88hJzXORFNXoexMelmTW1VW0VWNO06GKI1/ezcftGjsmuXbt27fp6tAPoXbt27XoNdNB6x+X7tdnx4YNfvTejTQlLSiZNVHpLLndzQKI8z5QSJvacLGXizHnO+TDlmUr0JwxMKbYuSICM0KrXFRzr/f39y7sXn794eb+sAvPtD//s//vF//y//G8fffSRIyCjq9sZXTgAlJzeuL364Vvfn0v5f//8z9//8KO7hyMnl+Z1FXMnopKzmkbJP0DPeoZodNadzuc/BU9LKUWbOzMREVVNKSWOtjZSawOAaLa2tVB7eHhYltXMAAF8MJbfnLWc4ymCmW/+6I4WI+wWO6vtRMdHfIEH5B0wNtybmz90GJmDsm1k7AwBA/9uVuLB7c4O6C2qI5B8X7NO5C743lirS/cTAMQEw+PN3Yhd3yJzMzcCwIDgkR9yQcAdogPS8DsPKh8LMlV3j7CRSJCIyIvINTYzEwWAnHP82lpDxFKKg6ta2LKYIjz5jLrNjJjHXaiaCTiklMrkAKCqS61RaDzP0zALp3hhZkZANR2YHAiRjidkAgQ9La01VQVYkKJrHolqrZWZc0rTNNXWVDWaDYqImhFRzvn08gjuV1eHANyqSkSZ+/uKCBERK6e0/eruaoZI4LiZzlLiJtJqm6aJiGxtTQURr+YDupvpuq6AkJilCSFNpax1bSKIOE2QAcPEDeAzEgAs6yJihChA7t5aa21NzIZ9BWqtOeecUwRcRFQoIaWEIs3UACGnxAwqEqdtTkzuoBDzEzn3zaQelNGR5kVahp/dzXEWDj94UGP3MHnjY5c/jCkDH1eDMS0CTiPqPgi+DY2zu487ZlRtG3vZFerXhtHtcbdD79r17ZW7q9a6RsATuEtrIgaq7gYI0hgAQaojAScQQQTMxaW6KMD4dE/ZAVwacNoqnRAJehNXAFNAQEqX85Hu5qaROkXMbhqVcwBAl+sIYAArwGfH07/4q3ehvuFvXiU5JcKcylTyXPJU8lxKTowAKaV5nr73vTdLSjELzUwlc3zhQgBVUVVKHFPUqmoeIVHMxABgDmJexU94xfP00cMJra7E77zzd9955x9+M0dm165du3b9jtoB9K5du3Z92/WX/9N/d6960PuSOBMkMNrQJ3EEJEcSLhKmUubDAVNCJkwMyECJ0oGA0VHFXBTAzVSl1tODtlWk1tPRmhDgcjrVZdVmOU3lcK2pvLg//urd9x6OizuAbVRwYAyH6+vrP/7xT773xpuE9Oyzz5elIlJgx3lO5oGXlYlzykgIDmqGKIBAKeL/TFH6PRNhxNN2QyizO6eUVQ17ZDCVknKaAAAJmUlaq+t6PJ3qsphsdphIKP4tGcvGaLZkggGn+y9b2GKPeb4wSw9DcGfRPoIsYMRkRHACjrjn0ajNL3YuXMDns1m1AzkYzufLOIFLe/PZFbrFSD8yc+O2/OF8CqOvd3Ifmc1hjKXNxerbEs8W67PxGQC4lHC/XiYsq9mGx03dbXPIwiEfgic6eEo97BsRNci1+zxNgFBrDYe+mUkDUc8pE2FEQufMZbqJSQgiIgSmaUPesYszpi24YcuOQMRSUpkiSdkiHxociDFnHhQdCyZ3JmJyJMacEiCaGdIMDswEHEC27yMRYeZSSjSGQgBOiVNSVQQsxFu6Mo5c6ZTzVCaO5ptEtVV3n0oBiDMFiTClZKLgEFDg4M5MgGjgRJQSl1LC3VxymUqPi3Z3IpxKZqaI4EAzIs4ppb4hqqpxFIg4pRShGtEaUYhyGMkjVuZizqNPfPTRjoAUmaTDQz1qtQNHW8BjYg4AjWqq6qPAeouriUaewMNeP1LIexXBlsChIiJNRETEVaNCIjzazOQm2qqqRFT0vylb4zuBYUdlA0JMoQ3v+ndi43fter2EqGYvX97dUrq6vr59+jTlbAbRefccPqQa33LADdyByDRF9QwGMo7UDJ+IOH6M/n4ikSWNCGDualGmBhFpFd8PcUwHOgJCVnCVV2vLHIAQxOzz+9qMynzIiuSGDmq+NlHR5bQQOLgxcyn5/u4lM7lZYppLvrqag3QzYxNp0qZ5LlOZyhSfSYQURUXxKZOZmZiI3+Kbu6bL0h6uSmr1mz9Eu3bt2rXrt9MOoHft2rXr266GdKNy5DxNExNO08wETEjhK0HklCglSgmZUs7zPCPhwMUIyOYubdWlttaCy6iKtCbrSVo1qbVWNyOkWqsblDLNT96g6ebTB3t2d3r/k+dr0x418VhE8Mbtkz/5W3/rMM9ra020lInzQZoxlZInMxMVFU05MafgrFHab+4Gm+c3gggxpRSAMvywOed+jyRbS/fNhdN59Ol4lFrXZW2t9cbu3Xj5r6crX1qeP+AxjG6D2FMu4MKRfBEGcGbNF1guSmK7fODfuJ/DDqC7nfNyOReu321F6MyVR2DHhTf68uEL2P7Iyn1uXu+XnHprmdhTVcYWwiiKBYs9sFXnnhsPXiRxwNYByZ2Zw8/ere3EEJ34ABCRibaphVA/1uaDMPb/erNCtXmeAikSEUIEU2IynkpBBDUDd2LKufRoCTdw9gxECN4b1gXYNFU1ZYoYdFRTJMwpM5MDSBMJ+1XcgSP0d/RtFGG47EvOAKiqYyqg74mUspuraBz6nLKomukGC4wZkZjTRmnD2NV3CHj37zInJjPLOcdUTSKKJGhPNgYuAgIhmruYujkTTaWIqrE5ZGYmGuXVPkzsBKYYHZ96ODOAEyVOMQQjPPRytoOGT01Nw/vfh13Y3gnpDKDRwU3d3NwsMjbM3KLxFTkiIkEPV3F04GFSxtHEk2ibEtlmSsasibtDv2xodOWqtbZapVVV3bJfIhU8jr2KjFH6CoP+7kLXUYoB6GCIF5ebXbt2/VvTFyoSUNXv7x8O1zdTma5vrpFoXVbwdFFNdQ7B6pOdGB9MkFL/ojVKoICIcWQhuTuxQDT4jWndMVcaOV3YrwweXNvdIdFq7mrjLR8VwYn6/UmqOiW+nq/I1WNSE4BGlQ2CmWu15lIBwc2YqeR8PMXMKyXmKrW2Ns3zfJjneU4REkcppjERkSmllHOmjHQ1T4d5xvs6nx7M+Bs5Srt27dq162vQDqB37dq169suIWrAYkBlIoarN99EcCJMKSMiMU3TRKVAKcFqEAxErLbleApv4+m0nB6Oy/1dq1VbDYjjbgjAnHIuc54oZWCeAYjz4epmevJ0hfz8+a8/fHH65KUAAxOI9FVC6pEUKcH3v/f0P/z3/wMVefny5ZMnT56+OQGlF5+/nPJ0e3PbWgt/TcopbpCiw1rJpbZ6fzy6GSc+zIfj8SQih8Occ0bE4+mEiPNUAFDVlrWWnFMPNBjrj5hS/hxheXjQ1kytZxWfLct/HWHBR1hqhNOGDRPgDJ+h25Xjj3SJliN/oAMdukTTRJfhGJ3VdVAXGHgLOqb+9MsVg9HaDSAaFXr3OV0EfGzrO+5dewrC6CYHA6GfndCOAI/eqy/2vFwAGIHd5397ZkKkWA83OI1iXARwIuh2aRw4EgZK7Bu4/QpbKkhnkb4FswzbO+R8UFVpjRMz0ZSzeU9mmUoOt1TswOj4h0jAZIlHmgRu5s6UUsQ1iIgZT1OJboHR8DDnTGFnNgMnRjwcDgggIpwSXoBmHOZbQGQinkpkaDBzrVVEppJcXdx5ukJEc59LBgD13hgqpZl65CVGiHnJhVOKeBl3zyWHGRydwSnlFFMvrca9d5B4jNkNB1dRJJywlMSq6qZX00RMGha5iPF2c3dCilkfSkxEOWU1FWmqlphzyWaw5d4wEwCYqpqXnHocCri7E4/zpMe2ODGNoeTDmt/Hp7ubuqqNw0pk6BRnKMX4SJS2evDzVMw58QXGWebuLtLEzNzVNgC9SmtmCm5wfvc4t3FLjj+fVuAXP/91v/6NVUxI0dYLdRyyv+GbvWvXt1v4JdcgNINlWaUJJ746XKno8vCQUuKUkNBGLlEUzazrGlfvmINPzAA9zQwusPL4PmAxrx9fdZg559wrS1QBeudbMxOpHJcLBxdzVVMdoc0Q5V3uLgrVYF3FTG+f3MwMbo3c0aNFsiMAE5mKqRpATCTGFPLd8RSOZmRsrdXWeGnp/pRzJqLEKeW0lcNkzvM0397e5quSCmdKAEZ3SFm/4UO2a9euXbt+a+0AeteuXbu+7TIkYczANzdPZhSUXkZNzJsXVluTuoqqqpgKqFlr62mJtm/LsqzLKnUlcCaccqKphNsy5ZJSQU6cS5om4IS5pGnicrXcrb/4q/fe/fBjBUjECACiQVq939jQk+v5+9978wc/fOvX7773/vsfvLx7oNQQ0/F41KzoGBm7YXcFxFZr2EuZWExbaw6OjVptARNFarh1WqtmdofInACgNQ2DKECHZXFTRYgPd/en0ymQ9DD8/k5QJVyUgzMPVDpIM2CEElCwOTj/ES9ecs7cwBGxgRvrxc03/UUf9jA0By46e877e52fGC/uNmcIK/Pwbo8XjLfucBrczLcsjbGYWI9zQT52+uxx4xne2PGSDrI3Q/jm4wbY7hM3do+ImIjPhlbvpf9hVY176C1kuj8SaR5EmDPiCJQ2s86yY9Ex95C27WBORKhm8d4iLZoQRnZHpILELToiMQMTAQATh5XYUy7j7eLdoaeRcOB7HHs1go9LSrU2d2PEzIkAExEgMKKbIXYrsYOTIQDjGMZmCkCRQpITMxMCZx4ENnIqEIPtppSJ8BRvisCJHUBEckrM5Ezm5uZ5nlW1tTqVzInVLM6FNEXWtqsIAHGaYjghIKecU4pk6tRXzEU0MUcqiAIiagxxc6dw7RO7W5+HgDH6Ru/K7djFxEpUdCOgURjkx0TJaGS1TUcgGozxY+7bbzGQAlW4mVuADHYyI0EwNzVTd+sAOpbtlwP+FeGXXRm+QwDWAcwBwBMiARicp2o2fWlhyK5du745Rd6ZQl3X48MDIpZSbm5u+oTo+PSlC0WABjMjIjEhoI8+w6Ox8/axj3wxDx0fcEToozMBIjITIpgRIblba01tpPjEInr3WUAgdxC3l8fTZy8efvyDN9Kc2VMCZyQGQiBGSolNRbW5g0FvbguAyGzj+0gqkkT6xpupWmuCK0bLABGZynQ1X51ORyovYLpZPbO0RAXF//v/4u/8l//DP/5Gj9GuXbt27fqttAPoXbt27fpW62c/e0dNZi3lZppyKm4EDG4ABq4O4OZStUqrtdbWpEkTcTNX0yaRwVpVzNTRU87TNF1Ncy4l55xyYc7I2d0plXI4OLMzO7Ea3x9f/MXP/9V7H3yIhEjsDoADQDuAAzHdPnnyxhtPb57cvLx7+eFHH714eQeYAKku68prXWrtANpSSgBYWyUkYtpQULCpuK0xt4jKRSKz6EkjKWUiMoPwnybmsOowETiY2d3d3fF4ig54scjfaY93VDwUdHSYeQHBz8R1+IRh4OQtrQK2R8PN7JdRzOOh8X7hd44OhxcpG48K5DviHb0Vx7/jLrCHrVxuh1+s40azezJC35djuehhtQ7QPMzcW9i098ME3UkNw2aKCECwNTf04Y3adgEi4ADNW860uaPDyO7ozw2PuG0Vu4jMHNkeiOidzgISAIJKJ2mRIG1mSMSJ0TyIu5k79CjM8Cw7AKrGoWVEohyhDm7uDom74g6fiFQNHHJiNYu+i4O1K0XrTMTYn0zjbQiIWBsgQkoMCOFTYyZOiZBU1Q1i6ogDEyCmnkuBZgrRSW8cmJwTE2lukQTNROauGGg32jSBgZaS1QjAOFEEbMSxTokjt8TUiCj6KJqZmxFzTAJtY2tEhnbDc5Dwfkz9PMxhw7roANCH0vDjufs2wYJAhA4ECAQQdmy3yyHS0WfkQ8djPlJTtgE0JnAGuiYiZwo+AuDu2ieczv9ur9zO511nmTsgxnlCl9j+Qvsu27Xr36ri49Lqst6/vLt+cpMSp5xEpEmLwH1EBMJodRy1Lojq23cg334EAIwCou3Bi+axI1YLzl854muYmbmpIZjq+Ba3XSfOZVcA6Ajq8Nn98t5n93/0h5ITz+hEmIiZc6KUmEviaHJMPR3OzAwQKSU1jSI5NW2qamoagViq4wPLTKWtjCCJT8d7xwfPR5tuuUmamY31sops165du3Z9i7UD6F27du36Vuug1y/50z+gn95ezbac1vUuWQVtrqKm6qZmoiKqKmYOoiZiouLuKeVcpjRN1zkBsSOmlKZSDvNVVG4yZxxID4igZF0Wfagi9vyh/qtfvP/P/9k///D9j4gSGLlZAF8cuQ+M9PT29vrqSlVf3t09f/58WZp6c8fWGmNblmYj8jYxhbW5WjVz5iB0tiwLEV1f39R1bdKIiDkxk6k5AHJWB1UHx7hLAUBVba2hg6rWWo/H07Kul/X2v51GXPOrhfs+imT9As2cDcHBps2i0hV6fiIOdyd2W7JhT61wjHs2RPRhlfZhI8Xhpx7v0tdsEGbHM33GjVcP2jtW3MeKAEZmhndOaMEBYQDt/kbDgoRwiRpxW1R/j0GgwaOJHwCAWbe0ullP3uhhIYBE5IjWC3tzLnFLa2bO4AiqBu5IYI5oQEQREb1lVqpp8E93cx9TA+RqLqZqK6cESKoCIGqOCLF8TgmRxCLaEjklN1cHEUU0Zsq5gPnaTq01cJimAmCqzkwIZBC9E2maZq+1aQVwcgzMDQBNDYkJsIl1cm0aUyBTKQggqkQUd9pMKeVk5qbeVIhSSnme53gJBPJFgN5lsaacmRMhxo24E5Zccs61NXK/LiVqq1trwbLVzQE4JVVTN0JMOQ8beM+ARsSAv0gISAZuqohoZiLNzSKfWlXFg+xj7EwAQMLOLkTjcXfpoyZ8bH2cupmfiwLOJDqQObiZe7Qd3LLfYzrG4cKs7xvnwMFHw9e8+ejPp6ePiRsH9McQ1cdwvkTn28nznZY7qAL27qL+ilf8d60f2bVr19cgB4da17u7u6uba1H99LNP67KIKnKK6dCU4vvbOQM6/k2JAcBHCFFUsWwIenuDUXODAKAi4M45x6+n42LaTFtKBRG1yZgJfnR1CEu0OrjDhy8bwP3NzUc/us1Pk93kdD3NV4frueSSU2IsOc1TKXP0bxBmBnARIc7dcB3fDjx6QEiQ5/A+9y+0xInTulQxNODGIAzuXhPwfs3atWvXrtdEO4DetWvXrm+1SPl7+nYqfkhJT3dyuncXl6ZSRZqYqpmaBp0jToVT4ayWAXE6HPI0US40ZUwZmNGROZVpCou0qHYLoam72en+eHdXT6savvfxi7/4F7/86MNnp2Nlyhod1WAYdREQIKf0Rz/+8RtPn3762bPPn784nlam4k6i5h494iR8OuhoDm6GFHzS1awjUQcANDM1UzVEipiIR0zEIZ4LESlg0bcdVa2JNmmi4l8bNrm4STMAClh2acsEs7gbO1tD+81feJQxQpO7MzlSk5Hw8TZ1dAZobsNa/AUADf0tu2MROqcDx75Om+V78ynj5TPHXMEISLANpsd/wwP1ZXth/B9HmoEPF2sHzNA7CvYnD4w4qGO3LIf5FQFFNG4uAQEFsQ7MSL3yl4bxWtUQMaIzAIBqj+ag7hoGkd5tMveWgDLKkDG61DFzH1QqUb/sIxAzlFJ199aaivZVNzP3UgogqqmZMTMRr+vaWh2Z3dhd10SRGAMAZNrReUgdEdzPCRLeRM02SxcRqHkTeWxS68fIzMScSGAMO1Eh5iQqIh5ly4je8zp9O4iwGYARc8pEuCzL2Uhu7qfT1iVSVd08MatZkwYORJQ4xxZ0Szpt8x/D/z6Mzue389Hscxtl1kf+1lmQCAnJ48xV688IPN1bbOI2xKMjZZ9qgAsfc5//cADQ1lqPfu7JM32W5AtseSzhFQb9XZe7Kxh52N1hB867dn071Vo7HY/SJOf09Pb2s9a01szZNOwHfcK7f5Q4RGMPTQmi1sENkYj54vN/u47GF5Q+E711b95KrQCg9yQAYGZHjJq78ZVhfAr0GDA4ib9Y5NO7ep1oOiBqk6qnU0tMTMAIKdGU0+FqTomJMedMhACeEidmZjI36814MZfO1r3PcLqIIjgCTrmYoUE2mq9nfu9YjYgZ/8E7f/c/e+cffsMHaNeuXbt2fVXtAHrXrl27vr362c/ewZVMDVJjbe101OXkoCai0lqrMiyIyJw4lTzlMuVpMgfidLi6osRABMyYEqRkVdwB3bTVttbWqqq6GhOatLocX7y4W1ahfPWrX7/7lz//xcuXR1XETGYtfKydNxEQ4GEqf/LTn7759On773/w4uW9GhxursVwbQIG7h7dbEZcQLhbgJmJRvs4w8NhDrsrE0HOkdQRTs3AskQEDqrakw8IyZGZ3dHMMRqsmX45Rv3q6pkQG3+1wXxjTbbnBCwGgGFQ9lcXcwGRg0g6bvEUZxOz9TLYDbpHifzFK+FMiPrdYqd8HS73N+yLALxk0Gd818cJdURMvm2ov7LNQVp9hPQibnCx3+XiiJ7eoOuIUekwssPFsVoddDnYVv/rbqZx3AEhjE5IxESI0Fqzs5MLvTvfIQYJETUJ/ugRzwL9rpUA0dTMdCsuVlVAnEXCAsbM3Qo2wi7jX1OLZoDTYYZoQsjMzLW21pqajqBkM1NOaTrMx+NJVUvJ0CA2ys3NbNEVETil4QGm1sTMWhNA4JwI3azW2qKB1LYasXcRAaC5u5qWlBPxWtctAcTMmrSc0rYhQbXDCh0H0dwjgXpZ1pQ452KmItJay7nEC0XEVHunKVUmJiLCOiBy5xOcyAFMdfSudFM1szGrsZVin7NnzNxt6zJIvUkWEfSpI90ABlF4xHEbT9tMB2w+6m3ep0ezDENca52/4/bys2m6j+KLJJ1x0vYR+fj0vPD4f2fk0I3u7ts1adeuXd8uqei6rm1dr68OP/qDP6jrKiLTVFqtVSUm38wsvie4u6tGztGoVTJmIuZ+GaRXp+BGkwnvoUzM25cc4JgzDwCNatYQXJuj46OLhQOCAShAczg2FMi5FJfTWuvptJiom6IruBLBPM/zXKa5pJRLzmXKiSkxJU4GZmgl52maDoeplERE5l5yJqJaq6khOE2MwOAEPNd0ePHhMxEpT250Fdi1a9euXd967QB6165du769Su1wPz2/Pb7VpN2//FyXO2+1uQESpJmmw4GHe4QTMTNlTplLaXUFN5oP6AYiIGbHRaWejsdaq3m0Ite11taaiKSckdDdVKzMhzd+8AfyL9//8NmzxURQ1VZDBQIwAAAESAZXc3rr9uqtN98A53ff/Tjl6x+8fZivr5t6rSK1MXPKWVpDxDJNrdXWqjTJOZeSo8lMdFdzBzNlTsycOImqNCGiCI4gQjNvrbk7IKSUIi6wrvLwcNRWg0sbwBfKx7+YZYpf9mv/17tjuCc9nGv+x3O924q/sFR3j1iBgNK0VfqHSRkB3MA9TEYRJL3xXt8WAIg4PEqXNiXEM012AHBzdRstDaHbRH14kXuXIt8W/kgGhta3xh9tiXUDqyHShWl0C+i+8Jf2vdBh5eWWOIB3o7FFXa17z12IrTMz8YaIRNFaDtQ0ej66m4gCOP7/7L1NrCRZliZ0fu41c3//8ZuREZFZWf9V6umu7un/btRiRgwMixYbphcgVqDeAEvYsKk9ICHYtYRYsOteIISE0CwoJBgEIxqhZmborqquyr/IiHgvIt6vu5vZveccFudec/cXkVlZWdVZUdX2KfPFe+7m165du2bm9zvf+Q5RADTPLHbHjsCEpCagquZV7RAAxHXNBgHRDPquQwBiRiQRSUMKMRBRPyQXaxOJW593fZ9SUtUYY+AAYKImYl0/IBEYpJzMeqeECckATS1LVlESVcSuH1zR7Av6GIOp5ZxLTGBIgX397OblZgaqpn32EpcqiiII6GYd7mzuSQHMBIimKlkRUCRn1awaQ0AAETVAVktIroUxAAAgAElEQVQ5O5nrJDubZRFDjBxWXa9mTJxEk3Rewc8Muq6HUmAKAakfEpTajyCiYgKA5pkKiESoQ0lGQCwmMYXc3xDejzGYepWMsQevamVm6t6kGzo9N48WgLQmmOul5PI6b9D9sMss8oxsU1MxVQBDQmZWQFWx6sZRyWUscnzAGu/ZZKhfvoZ/LPwisLXm2QjXgk/XrUw+zUD9tLaZMOF1wKe8uj/llP7RrdlLv2z8qqayWFzNZu18fuPg4MAAVDXGsLO3F0KjakNK/l2DiEzFTJHIE8qgWht5ZQG1kmZkNZ2ppLSYjeE68EAvMwJRiYp6yQhAIMqsG4k7aDDa7htAynp2fjUczXZmBzRkjsjMJqqSU0oIQIREoIBdn2XZew4TIhBSCAG5SLKbJs7ns7293aZtESBECYGJKFAk5siBkRkJOMzanbtdvzq97C97CJMP9IQJEyb8HGAioCdMmDDh9UWEEFc3CaUJ7dBdRgJqo5khNxgix8jEgSkwF2sLQERSAzWVnGW5tDTY0KOYppSHrlutUk4GykxAkFN2JSkFDNRwbJp5g81+M98/verffXTcpUFRxS1WS148Oj12tL/31pv39vd2F116enJqHGIzDyECKgAEYuYQYhgQAYCZAQKiEWIIIYQACFaqy4ipYQixaUIIiIhDMgMuld7QBavMOFooEFIE1qyEvvD5BPHzj1wlVnYVq71FURZvizBx5IHrZ67rJtd9MC3ezoCFJ3X21U0pDLQwdLjZP6zczwYX5+SvFW58vTEiITnZPZJpVUULW8vYtWnHWue8lkVv+BuYeXwB6WUjg3Vrmym6lROnsbGyl+oh7IXyygJ48wyJCoARIjP7n8XegsgZxhjD6DLhjKVruFRLgcqmCL4US3+NmBHQ9drEjAju49E0DTGpE8VmvuJtmgaJYowiEkNkZkLQRtVdxhGd5xUVVSEk5hCbqKqUyYrvCsYYQwgheHazx0WMiF1t6y7nRIgl6IAiriumEiCI5fRhzoReldAl21p/V48JELdsyipMhEgRIDCXk4jFjsPPPIWACEycMpJZ27aqmlPGQAhISFmygjEREyNiyhkMyBOhiya2zAaf8iWm4VPPTE1LFKSaxqwJ6BoOISJ0d+H11CszoIjSR0Z7JDJqIMVPUGn92hWH6FkXBgSEYArAfvfIOecMuq6/NfpKbJKqFeWC+UVgkH9yXE/bAADYIOt/DNZ44pcn/CLhR94fXhmI/gztfMJ29W6s0q9WQ98TUtu0s7bt+i5wDKEhYjHjGFQ8tYjNxMAIUUUki9+GVZWoGmyQB8XXBDS86j5AAAg2Vkr2iDgKaU6qCqbX+4lgBln1atmlrO1s1jbWkjVN9GIlJX+uaK4NAIZhUNVSDhFAvJ4tGhiIWM7aDzlwAARmjiHEJkQO7tcROcQQOTAZztomIF0aZE3f/vY/+va3/+xTjvmECRMmTPiZYCKgJ0yYMOH1RWvzwDZr484s5ovz+e5u00QEgDjD0BBHzclyZkZVk5TdIkA0S0o5DV3fp77LXR/UQNQ0u4EvR0aMzCFEagPHpmnns3Y+b9oWm90e2hcL+/DJ2fd++GSpGzJdBEBgIgIysdu3b3/1K19q29nJ6dXp+WWc7cQZipm4JTWgiLpVq6ouVyuvtaZmMvT90McYEVBVV8sODXZ2dkRMLaeUhmFIKTNTiCFGHrpeRWOMZioiw5CIOHDoumXXd1mS12Is8uzPgCJ6HonmqireEAQVtg/Q7a9HuWdxqXAOzXwZZlAHTSt5TJVLkzKO6/YLw1335XYlYNXlGdd9KT1BBERiAlhThLAhQR2JZn+RqCyVSwUis2INQeQHUsoT2sjNoVpW0yqi3mToR66wCJbRjVNeHlFf55YOkGf6i2oIgZkAIOckOYcYyYXQpogYm8ajESEG9/fwxgix6l8VkZgoVovnUfitagDAvAeuqzZz32P3loCi1jYwIEJm3tvbAdebl7gN+GZuxFGFYe4uAkTUOJmbs4uaU0p7vMPExOTOECWCsTbT0LEAVAiRmb3Y5mw26/pBzTzWAq5oNgOAGCMAiGQo8nKVnM0s1sJQWTIAhg3zDSDyA1SRlFIstQdzFgGA+XyeU+q6rmRJMEvNO3B7a3fF8VF1TXzViePaiMNn/abfs5kb7Fi1hobqN45+4pHWs3EtNy52zZusRyWgfbaUKegMRW13nXJQig36Tz+/knNOfd+PJTbXl2PZ+6chgP5Wk9HX1M4TNz9hwuuB8uXC1NIwpGEw1fHhTohMZAZMHGIY+qRqnssCoH4/9QD+eLNFxBCCwfr2+2raew0FFSJCImRCIpGch0FFVMms+Fytb+4AYrrq+ywa29lhO9ttqG04DUP9/mZjsURmzjnlnHLO3kl/bKkq1T/PFmcpJRUldjlD4FJRwGKM8/m8aZv54S2e3dCcweB8H2erSQQ9YcKECa87JgJ6woQJE15T/OV//18LqgU8un3YIAywjLOWmEQUzCALGMjQydALqKQ0dB2YquQsue+HnHOpgWaaADEQ006IDceG26ZpZ6FpADE0sZnNuG05MjEiz85OLv63P/9nf/XeR1eDWZXqjspaVSWwiHbn1s23Hr69WCxPTp5dXF22BqFYBXi19ZGOAmeNYwwcGACyZLc+ILdvFkPAPiUgUrOcU1lnIQAYoqEBIcUQnHcbhsEJ2eVqtVwul8tlzvknYU0quUyVWSViKvXRtthhHCXAlU/eUmiOzPRIFW+8hUXOTYi12N6oJ95odWy6ijm3bUDGjFk1rcx02WF5ox4SbnXBKke+ZroLVVozbguB7iLW9Qa49umwUdAK6+PHzZ5dk3Ovtd/elFPr3hcmohjQCXAwV7ubCIIhoRs0wFiS0cloUwRDUHcgcbY0BCZcV3qMhOaulohGo0a4dN8rMBZrj5yRkDn42Km46wQyAIClnP1z46nSNCDRLEYizCKWMwMwYQzBLzkRIeIYokv7s2RmRoCUc2QKgcUtboaBQQNjCJhTUtVZ26iCiDB6eMINUpCZpVxu3n2YhViLcSqDMZMhApikhACzxu2wgZgDEQAwADJh23rUAUwjMzANQ0Iz2BCeF9kyuDO7ESEYGJU6in5EVbkMAGutdLV8QQQgImJCoso1X1PS4pp13jYWr7N9MxO9/LdpBVMJaP/VAEwlcAjVBtokg6oUf5jamPcXAWMMO/M2MoJJzjmGhgK5Q/fJ6aXVCMzfVkzM84QJrw9q0A0AwIah77pV16887rZYLIg4xD6LIRHHkJMYlIeRmvjnyZXONeiHiP4lSrSENmvJgXU4feNLjN/03XMNzcPiqh7l84i1Pz38zlkSYwxX2Y7PL3/44UfD0c7RTjOLxAiBPGcotLMZMxITEnjOUc6ZCAFBcvZwLxp66DelLKIqNpLmHhPOOUmWy/NzDA0tVZvuIvOKmiOb9VE+9zM1YcKECRN+PEwE9IQJEya8pshkYUV6hPt7u5A7GBpkErMkWUVMB0aSYZX7JZnkoR+6jsFcJpxzFoMQG2bmEAyZQxubWZjthHbGTRuaNsQWXWXcNMasoCkPIvjkxcX/8ed/8YMPHw8GPHJ2a0bJEHHeNndu3rr3xps//OD95y9erPreQkM5D33nDKOIjTVtcpa+79tZG2IAgJSySI6xKF8YAwIaqNUaa65yHWWsgYiJ05AAQFUlZwAAxGEYhmHo+17lJ1h1VD0wIOLoAk04FuvDUR09GnGMOuVRDQxbBPIWlzxSz4XoI3dYXuuoy0pzU+AMUMWbax53Q5okqpZt7F95W10mbCNzjrTRXKX0nN0eV52jk0YloMGcKiaAaq5RycQ1U4jbFPNopHBtYEfCkWBkG8tAVvmsOoeuVuoz+rjmXJTiVF0oVRXM0KsX+urX2XGBuoZGQgBTUANTL2+npn5co/zZZw7UwobFE9PARBTWnaOiw137QIiqewkjMIF5FUVQIQiqqjmV1bypj2kgV/wbmoEqqBKAqIoln1qgWbyUYhPQFFRMytVbTyu7eF2rJpqaBgAHSVYdw50KEDfxIATXjJv6bAZVPxYt25XQghVZN/opxvqfD6IzCmWyU5nENjK6PgtGC5lKCPv05sBjUKJ6X9ch34pWQB0eK6RG4X9tnKKjILpOrCKHL7J8M7BCT3MIIWdhLpNknIG1xwjYNvE3f/kb/+a//jvf+tLNfHn8/rs/+PrXv3nnrS+0871//t33/43/4D93O+y/zajDvv4bYCKlJ0z4GcPlwF3XLZcLYm6aBhCziNqQxQwR0yBiCKgxqoqoGBgjBSId769gRCSSwUBU05DGMrzj9xCE+j2oFhBex/rANzGya7cJ72ENMRoksRcXi/c+OmY5yv1sxtBGaiNH5tmstbaNTQiGxEiEMWAMwcPPALE8SID8q4NbfZiXny25Oioi/dB3fd/1XTYYhiHJSuOBGWTNsLJv//EffvtP/ofP7/RMmDBhwoQfExMBPWHChAmvKRSljxSd6NRkOQ1pEMnDMAxJJSsZ5KGToSMTk6yS2xCJCYl3dmcUIhIjBwpNaGexnTftHNuWQgMYkBmIgAgNTDR3fd+tlsvLRa9//Vff/7//n794/PQpEug1FggAAWLko6PDW7dvHR4dXv6Lq/OLCyT0gmySs9deE8lE5J4AzpQ1sWFmVQFmRmSqVddAvUQOMhuwgSIiM5sBIQZiq06vzlqWQu2IZjb0veZUEkE/E1eCVQu85l+KGa4CunUDjHRt1QYVOrmSvJXuLYRd5ZlH0hnX74xmGiOqJUFZKFZqe/3u1q6JcENbXjjxciDrf0eS3O19y3QahdCuFy7+jqjj6R2J2pGSNABAp2INoHp4aLFhMPFugGElJquLh2ujoBhnBCYzyDkRBWImIsk55yHGyMzM1HWdqs7ncwACsKHvETHEUOZHWSpDJHKLFwRgohDCMPRmxtVVfBiS97aJjZn1Q8/sMY/kY2hmIYQYY4xRVbuu8w4hoWbNOQNCDLFpm5xylpxz9vxfDpxzXq1WbpSRs1ipyAd936WU2rYVk5xWpsrMbdt2q1XOOYSgIn5EAOAlE7MAQPYpbYsVAKgaYlI1VWGv3qjGIRBR3/eemOzndRgGqk25SNgAFXLOiZkBUERcjEzIWXJKA3Ox++j6XkTSkN2/GkD8tIpqnWQIACKCAEgIUqcasc9Kt1rG9Xwpc8azGWwsSGWmpWYgAACSXwg0Rm6cLFaztRepqoFWEb9LrdeXdKkk6L+Xsp7q4SjNbhziB0BVKj16yuB81r59784f/iu/+5vffLhHV6dXw9tv3//SV75w487dnNM7t5v/7N//1/6LP/0nf/3oxY9x4/hFxIbefMKECa8LzCCldHl5efvu3fnOTsp5teolS4s8SO6GwaXDkLPrm00NmdWtq1QlCzGZaUpCRGNSU/kWQyXE7g5LtTwsABigWYkWgwEQIseAQSHn8m2g+p7V3BgwgMtl9+hE9lq21EdJbYAmQBMohtDEEGJoYoxNaNumbeKsiRyYQ2hiICIAdMcqIi53/bX6AQFMTVNOWURUuyEvMyy1WYa946ulAK5ShzwxGxMmTJjwWmO6TU+YMGHCawrBDAYkYbi61MWL/vJMRUVykqxGZmgAJgnNgCiEOTHH0IbYcIwUIofAIbqal2cth8DEKtn6pampZBHJXmjNmback8rlys6enZ4cny+u+nWlGSwyGAQgg/ms/cLbD27cOMwi3TAg042bN0NszTANPRMhsUH1/10n2oPbT1RJ66joBUIk5thEAFssIYTQNI1kAQBCNjMVLWxdtTA2AMm5Sohrbv5nAZo5m61e6s8XYVX6WsS7G1QzIQGYoXqhNkD0yn1GWG2gi19FYQxtTY9Xgts2SwGWX5m5bFmHq8pQC2ft4+CEnZrptgAaRv6o/KjF70ZFKoyK1A2zDtuSQ48y5Y2+VjeU9U6KLtZq1cuqf16fAqtVB51TTIWuBTVFNQBQ1zEPCTH/0e9/YZfz1cVl3/ch0o0bN2PTppwvLy9XqyU2ex+dpR88Pn9+2cV2BuA+ksrEgcOQelVlYg5MSKqiZmAQwmBgOecqrNUttxQADsEdx4mQkZBQRCVnd2eezVoR8UwC1/EjkYdYQhKXpNURX3r8YFBTtZwVAZmJl6ucxU1C/HwxEQCamRTBb7G+sD67Z42XZFTJMQYCTCl7GcMhJSegVykTuqitOGmqqbowHEDVmMltwauUHj2sQSgAWIRwJYYAWcu835iaQBSQUP3MKpQZrs4E4KiAtzI1/aI2tNGVpSR9ywb7PMZiitO0b2Z1Io9z0bVvWObjxrStoZVNBbVfAqq5aOPMymfWzDgAIFhgunPj4Pf+7jd/6+986daudBerpokP7r+1d3iYUnf24vmwOv2Db729SPpn//Nf/Pm/+OBj7xMTJkyY8Lli/eBNKZ2dnd+4cXPWzpqmGfqULTNTQw0S5ZQBMMYoklVLDg0BEpE/rYgZAUTFy8+GwF41oUqeS+hxrPMMgAaqJv5wMTVP5fI0oxyDDQnMyySXoCMAKJgArJKdr1R51uzu7aIGTBE1MnhCjzs992lYrVZEiIYxxhBDLEURMDaxiU3TRObg4fvAHEIIMTJzwBDa6Fz5bpb9bCsJw/yQ2/jk9Iqbmcrf9lyWCRMmTHjNMRHQEyZMmPA64jvf+W+G1SKYoGB3fqaXp2l56UyLoSFFYkYiRkZmCiE0s9jOObQc29DMABGZQtOAqEqGGBRMs+TllfYryUPuuzT07kKraqIGIYbZbr8cri4XV1dDGgwQSymwSjuRAQPszmbvvPP2wcH+YrXshkQcbxwecWwNMPWDmRERx2BmIgpgRETEw9CZaRujC1GHYSh6yWomOJu1iMhoMTbtrB2GwdS8HrtqofzQXa1Vs8ji6krMkMj0M1pwbHlIoGHxinBnAEDU0TmgkM9ASIpKAIaoiM7LIRoigqJ5wTsDUyMyI0TForGuNBxuENBbWuqRMXR63m1tqZb4c4VoqRpnqoX+dvnS2vAWR0rZYLQGqRvgeLTFTteZR9wcijWXvzZehHIMRETOxbprI2gRKBXSr0yU6uZh5tpcpFp6iFxvq6qIQMhNgC/fnv27f++dN3fx+PHxs5NjiuHBwzcOjm6JwrPnz4+fPJL25j97PFgejl+cZTMXz6oWmXzRxUMa1eY+elSZ9yTiE7KqxVFEUs5+CDjabhTqXbMoM/U5Wy3052X+VBUIiWhQt6EsBjIiEkIIIaQ+pSwpSyAGBFV1zS+krKZghrUkVFZRNUCatW0IYSy+5OkCKqqgCDYMg6/5nUZHAEpCRCGElAZRjSGIqohwCAagZpireQxUU26ftqpmVmyuiYgwlWuzojppcDByixIArKI2BEC1opCrGvtKcVQH6NqMVXIZDBHMkxuK88zYnoEHIDY00/VCqxeGsxVWCeg1E4NuxKNmls2ySBYVdSbbqe3KkwMg4sHezte+9ODv//6vvXEYtbtEhNt37r714IGCPn92/PzkuO+7w4Mb/94f/ctxNrtcdN997+THu4lMmDBhwt8wUsr58qrv+t3dXU8yMzM1JQ7zOOuxN4BZ26SEqkxEHqALMSIAMyGSmaGgJ5A5AT3KAvwGvU42IiQkMcmSmf0LGDARIopm5EAhas62WfUZweOaAtAJLAbM3Mbdg4M5B+2C5UgIJuo1qlVFZEhJkqQhhRC9HHFxr4qxaWPbNjEEZkLCpolN28xnbdM0wT07mIioCTw3nCnBwV6cty8uFtb3gzZ//Md//Cd/8ic/oxM1YcKECRN+BCYCesKECRNeR/CQl/PdnYtnK7RWVpwSIjVN5BBCjIZoSMAUiJhDaFoKDXLEZmZAMiRVE0lDP+ShH/o+5yyaTQRzr7mX1EsawDQGjk3TzhoFanb292++cbL8cNGnpIDMgSnn5HpNRHD5IiHszNu333rYzNqTFy+Wq1VOYsgWDBGZKOcsIsiMiL7ycUhmMwghFBouC4B5cXM3QwCA2ISjeOSmyaCqau4kIVlVJMYYmyYw98NwdXnZ9X3f906EGehnFEE7cboht4RNdXJVYhYjaH+pGASjjTXSpJgMiFRrjEIsj50y99cttr1qUIwN3Cibmbl4UxRVeqHUi4ocqfgVqIoUArpsMJLXtZsjrQ9V3T26hjj9DaNJwVq65MUGt4hkLfaP1dSjUrxFlwRepGijLhy6xMlZySJyhqIZJ1/V+k69scD4xZvxP/mHD2830MT5wc3bi75Pw9XJyUd9zgc37ty6fdu61VVvX7w9//Wv3Xv04vLZwhQZCYvkFSnGxqBIexGpibHWNSJEAsJYSmKaO2n4cbulJHrdPJ+NKTNzjMFtLXwpbmBUHbyzqLcwRghGjb/TqExh7tyrnyUR5kCEIsqBA3NK2cyIUNTEzNTaSkBbrQblH3Y1WgjBT0/TNITEzKPTRAjsZ03BAMCl0yJKjIUJcIvk6gEKaqWrfm/hTTq4xBy85z4JreZcj34uZQMtYQ1C0rW+f5wCpqblGvItixUNmYKhYtHFG4BlyVZcojcusXL5ASJKdfioF2LZz2i+kVNKaUgp5ZRLAasxYuJXHEJgevv+3d/99V/6jV/7qr74cLm8nM9nRzdupW7VrS5fHD9erZY3b95+50tfofnOv/WHv0M6/Mf/5f+Ys3zmfIoJEyZM+BuAmUHX9V3Xxxhns1nO2g0DqgWMBqCq7rBUrJlETJSGoXzn8AB2luDmS2ae4gMARMRFfQz+dAOEwCymqdo6qRoxI4KomCoiARGQwqiYXqdUQTZYZD0+u7y9196cHQEwEzRNQCq5Yf44KYFXKdUsxvwrfzqkRQJQj2S6BVQTm6Zt2radtU3bNu2sbTggcjLmZsXcKmZLckI32nT2szlFEyZMmDDhU2AioCdMmDDhdQSDhauOYzuftSYLato4a0MIMTaxaQyw0L2IDOAEouYh55wl5653u4aUk1fqc42zmcZARGgcYtPGGJs2xqYJsQUKYb7f7t959Pwv//q9j1LOa5FsJWOc/Wka3t9tj24crvruB+99+Pj45HLRxXbH+mTOBTo313drVrS4xwoiDEPy9ZAXmiOmEKKqdF2Xco59ICJQMNWUEiAgszdpCkkyDwMS9l1/dXW1XC5TSpuc008BVgRBm1XYAIGKtHQzXRXW5tDjQVYBdSHKRu8SAwDTuhYUUURQIoZixaBmaGoKWswpYBx3VUPU0X+amVCx1mSrNo5Y3ToAvUJ9YRBdPUrrno9Wj2uhKG7szcZ/gQy3LBSImAtZXvpiLsIyHEnl+sNcp++15qri2zVWTvtaHr5wa+cPvnGLAZ4/PQ733jg4PKRAx8cfLK4WJ8+eDlneuv/2O1/40rvvf3g5LL94u/l7f/dr/8tfvHeVECh4g0zsevDiEIlIxE7/ksuQzZx1FcmEbotcPGGyZLBC3Toh7aGAqomHLNnMqE4ALQUSaSyHKJIBsGlizuJC6VFMraZOghOSVfp/1hSfZXdRAQAmRkJoYx32kW6FIqMvfD0SERNLrcTE7oGuxSylaLFVAzMguHcNlmW+qbmoeQQWnnrTWKVuuT59Nk5jWM9FcLPPEo7BLVuXQr2XWQm2npj1g+OctOoO7nGL6kxeTT6KiU1psQr517bO5spzyeMPD8vUilnrrt67c/Tbv/aN3/nlL8vFMcrw4P79nZ25pP758dPl8iIwP3zw8Pa9+3x4+Oy99x+/++5u0H/4O1/9x//0+/2QX31/+DkDfszrE8E+4dNgnCcfN5EmfF4wALDlcjmbz/f292azWUqSRACRmd2Zyp9iXiEDOJioWsl6ATBTEyIOITCXNDVmqFZQXi7CiWwziyGQCSAQMyKqeBYRkGH59pLZvPjzGLmu3cwAK7OzRXexXKV8gCqIwkxkgASExcasYUZAf1JXaLFWMqk1BMTTp8x0SH3Kw3K54BCIAxMzMlIwjrxQbfeHIWezg9W7qd37/M/PhAkTJkz4lJgI6AkTJkx47fCd73ybhz40ze7u0cFeqwtocDaLgZg5xBgbgEI9mmZLQ14u8zDknPrVahj6nJKvOFIaBneMDjOgoMzczJpZSyHs7u/Pd/c4BC9aiKFRmmfc+ct3n/zF//f9IQ3mylFdryv8585OPDicz2bNh4+P/+p733//0SNRPDyCbpVyFiPzVM2snoSPLskRkbZtmdlZpbooAgBgZjVNKRGWIuxuSw1gxMwx9v2AgLu7uznnlFLOOQ1Dt+qWy2XOyUQAf1rL48LneQ03K0xzLTdY+LRipABgbt8w6osBwUbSnerRlHaLHYKzndXheV2v0P2jK0PnK8EN8g5GRTWAu/3WunylnaqULm7WNpKTa/p4TUCjuYa7tAY6sn3O4Hmro5x0rKhYStsRja7BttG/TS9JK2QglaZGpwsDRAyBBfJOy4d7s8DWrS5enMCBymx378bNeyk/vbq6WFy8uNjZOdi/sX+wf75a7K0Wv/KFu4+eHb37vOuFgcivhGFIqkrOExuIqjPRTKSmQ84xNkwk7noB0DQREVVNJPuhqSiYBWaXRdfFOI0CMT9/vk527TPiuv7hbDZz/3R3BUHkENx8RkwNCV3jnFJu57Oya1v7h6hq0zQumt6KcJhJNT0nYn/RqiuIVykUdW9mEHFltIUQzCBT8lOWcwYwRAoxmNkwpHGqjJplAMB6rkfBsVYyeUtR7G4t41mukjVvyCd5jTgZ1vJWOHrOeBtYJg25YUbtQSWxy4wcNdlQfUbrvjwuVtw7QBVMQcRETbUw1TWvfN7wb//q13/vW195cHOWVxe3jvb3Dw8a5kW/ujg7BYSb9+/fuHOXkc7ee/fFR48R6f79h1/+Ym7+/IcD5J9/jhY/hjc0GE/Dq96YMKFic5JMU+NnDbPlYjGbzW7cOLIWhiENORtACIGZRXIaEtWUKi9j2/c9AITg9f1MCkONJYNqPKUGhbkGkOoHJSYpJwoEgCbm3y9EJXxE7osAACAASURBVOc89JA9MQu0Bg8BAAzBDBIAml12/eWy74akOiiImjIhEXAgQmQCt3qOMRL7VyAANEABUE8Xg6JU8EBj7rvVquu7rk/LVT9I1ycTMGCa7YaDVTi4tcqWxXA/zPruZ3J+JkyYMGHCp8FEQE+YMGHCa4eQ5qvm+VF+++jWraPdmbVImgjNs867vjNVE5Useejy0FlOklJOSSSpZM3Stm0TYyAO8wZDDM08zneb3T2ODYWAhGG+w7MW0VSyihLgYjUcn129//jk+MW5qDqdhLUIOVaZyxt333j74VuMtFwsL66ukEMMkZCZ1QCQEQBURSS7NmcUzPrvm4epZqKCQM7FwkiyEmGgSvZSExtn37A2KDmLiKlCpa9+EmzT19WgFgwI3ITADZfNnGE0rBLQ4kzh/sKEgLWiD2FZBlKhRglGGSdorcBYCWhm8uI+3hkVVUTdEC1j9fUtvJGSmUqhehGrnLWw0QpGpaktABTSsAhMR22rgYEWV14FMyAkKr4Zno9bjwsA1HzN6SSvgbnydOSfi/TbRi/p8jkzA3PbBjQ1MwmBZrN502YUurq8FIAj5N39mzcUmLBbXj598uFy0d28fff2jYN+WLFdfePB4VWXPzpLSUldQyvFZMJHwLXkrjA3ABNNNmREcutwsAxgYCJFe4uIOWUXfLmIeJSGbbK9ACDSAYxembYSiTES0XKxLONo7kScUiIAVFEcWWADAOj7wU+i86OqmtLgnpuqmnMKIfrvXvSwyP6dgq1ezz6S6gdY4gWm6n2ONT8afUygThlxF+l1HUaDjS2q+XJVGZtRsYzZICT9LkBuEI1UX9Niw1Iv1hL/gDGCUuYt4foKMDAFNfRpYtXJBeoFspVegPXKKP4dBn7Aqinx4D0WVdXqUF1k27M2fPWd+7/7q1//6sNbc1be3Tk4OmKibrlYLRdt286Pbu4f3NRBTp4fX548RsSjm7eXje3sPq+Bnp9HfMaev+Jj9nH89S8gNoi4T3hzE691eGKzx5+1o6/8HH78WxP+pmEA1vfdcrno+15ERUQlixUrZg+g+nbDMDBRICainPPVYtHE6FFVD+u5CNq3p6KhBgAgopSzimQRNR1yYiYAcAU0ERp6TJSIWJEMr3/78tuvKpxdrJ7tLi+X/V4wCkhqakYKUjymrOt6YgqREYAQiKhpQ9OEEDCE6Kw6IQGiKyE8qCuqQ5JhyF0/DH1OGYSitfPEuDy7ShTmYZ8w/6f/zr/6H/23//hzPT8TJkyYMOHTYSKgJ0yYMOG1QxCO+SZFmYfAMuSUJPdikovnaVKRnFPqh9R3OQ9UjF8VAZA4tKHd2W1nMyKmGDm23LTNbKfZ2XXnXhU3uRg0D6lfpb7n2f7pwj54fPn05MX51crLxFUyB5yjQgBEe+Pu3Qf3H6RhWK06EZvPd4mb2M4MOahyIDATVY4JEYjcN1DTkHZ25jHG0ccWEbNIX4TPFJvG1BAxbqik1yNSBZsaTCUDQEpJzRm6n5B+3vy3HK+aoSoCGWiV7W4TujAKjxHNEF21U2lYQiAuBhBOWfoYOvWrRW5cXJTJrGa/moGqqDpHtyb1SsNQFaFmpuqJtn7w6N68OHKCWvk/wtqvjWMeXUGgOgYXg2lVAAPGYDQq3w0BFcdjg7FTRGgAJQywrniIpbG1HwJaMZQAqEYhmjsDa+c7e0fBaFhdnS8XC4ovbu/t3bpzZ97wyRN9dnyyXA4HRwe3bx2ZpcX7T752796HJ+dPnl8uO6MQq1txMb1GRCZ2etY5RJeBF2Ja1cyGkMxMRb0n7s5hZr4Cd9G/m4S4LlhEiAkBU0oA4AJwFc0ptbMZEw0pYXWC9uUxIoEhgEvGSuDESeE6QiVe4EGUlMV3hDgYgIg0MSKS5AyVHciShyE5iVDPW6H4fTp4arU7tjOzn4KR84XqkFGcvNnZbRubGme3qtpaHIebl385lQiIqMWbxzb8TwiQmNGs2IdvGorg2Ei5BkqPALXQ6KabxLMnHlS+fmPuWpVJj5R1eXW9AYLFQLeO9v7gd771S19+cLgTGO3u3TeaNi7OX5yeHPdD9+b9B7t37w7nF88++PDk5Hg2b+4+fBj2bz7pTq8Wy9Fg/eccn40+3pwUn7KRT7mjn+Ko/hSa2mTOtm+OuLXVK4Tk9nF/Fov9V7S6/r3miFhNI4F1YKhGEW3U+39c3wGgppWUuxxSue1v7XijP1ss+ytO2ViSd9xu40CujcMvxgXyCfg0U/pzHgQEABFJQ8opIxEzZ5GUM2bx50LOWRABIOfMRIEDIoqIP7yQ0D2cDEw4qJqqmD9iig8G+rc1VRMAU005lae8KLlhFBhxrQZCVEvQrjMqDMGj7Fddvlilq5R32oYbRjREQ1CA+n3DhEwUBE0RAQnFgkgMgUIQCepqg8Ch1MuIoSFP9EL/SpkGSRkEcMCwFLiY8cKQEHa6wdqJ35gwYcKE1xTTDXrChAkTXjvEHEix4WSX56vV2eX5M0mD1x1EAFDJOaU09H3vkpbohcObHQ4xNG07n8/nu007w6YBDkgByCvEAQy9dn2/6lx22a8Wq+Xlql+F+dHzFTx6fHV2ej4M8lKPnKEyJnvjjTv37t27vLxarfq2mc/bHQoNEjdZACyUFQIIFJ4VCVNKq+Xq8PCwbdthGEQFDJg5ZVmuupQSB97b20tDArPdnR0AcPeD6goBoCoqiCSqy8VCRVPqVWXbB+KzwQrVVg7TCikLAN4HKELj0YUZ6k8cjZfXjY1kW3WRHrn7sgeXgBb2jIovMY1vWa1uB1U8XKnfuodSm817tN5hSVl1dWml+EfWfIPkgNEDuhLKhQ/UYvlNhIxAo21CVbEWn2dyPTcCEVrt8EhYAoyEsG3+4n/UwzDT4fLqIKvdefClbhYoUL+6GPrF8fEHD99+e//oMOckapfnpydP37//8K27b949v1zMRB4chu9yfv/8UrkhQrdnGFlvdxGuHBoCALt1JYCq1/fbJjPXtZM2zSZe8bLp5vumZrRY4Xiwnn1cIjZlfLCmJPvY0LYT8zhgCIDMSNj1fmnYrJ0BwGK5ZKIYAocwpNR1q7ZpmWis+rTuzUbPnLC+tqMiTBbx6EFg9gmlmwYaiIHJGYoyNXGTgF5P+42d2uZMo0rEV365zjMoaRTrox5JZSzT1cb5Um2tK01fpj4hlOEs9htehDDllCQXHfaIvZ326++8+Q9+71dvH7aBaW9/r5ntrJYXj588fXb8pJ3Nvv7Gm2Z6/NGjJx++F0J4+0u/tPPgwdXF4vz4+KMPP9RivTKyKj9HvNs25/9JG1x/tVL5mxzmy9zrT9Kx12j00K/X9Z9bsK3D/zSDYNfa3Oagt1pgRgRzTyAbs1Wg3O79UjL31fmYEasktXmmjakgQCDOWrJM6jZq6wvuOst+7aBwM0ECdIO53hwEqkf2Gp3KvwF8yjP++Q9CsTNSsVnbAFI+OVmtVsxMIQCSqko1g0oGZp0HwIk5qZiMz2HIMnjuCZRbdGJmJCppXkR9n0xFVcYQL2EGRFPhwBSiB7e1lH+A8W7pAycGg0FnsFTE+d5srw15IBACKVptU4TABMwl4AKgIrIYSgEDf6AwcxNiE4sgmpmaEA4OdnfaxmaRjBEZiVcpXSU9Ojr46GzxdCF6OMP08pfYCRMmTJjwWmAioCdMmDDh9cKf/umfDvpsRitNfHX2nLqz1HeqGUzAjAjYy69w0zTBnXBd48xNiwbEzM0scADAvuvFOjFzZWVOyVICETQDFTCXyyAT7+zMX/T96elp3/driWFZhBIiAhgH2p3N9g8PZzu7T54+y1nbdq4ckZhCMEQ3DTA1JGDEbJKyuIHwzs4OAOScobKQomJmMQYO7FXdmVnFPQcMEWMsdr2ecc+qhJiy805DVVL/lBaBZlA0qrimsio9uKFeG/WZ6w0qp7p+Caok2ClXvN7gmtfCscphUUlvKkex7rsSyONHrbxd2Vbc7Ffl7DeIpGsC6LGvm8S0m2YYQCkUROter7tcTIDHH4WA3hoWs7VMtWqtN3i80o7K4vLq9Oz89Pz0jVs35q09f6LPnh3nq0tJ6d79t27dfZMpDN3q8vLi2dPHt+/cffvhm997/8lbN5ov3dt7crp8dLoAQlWo03SLgizjg4Qbr5YCjBscnY4d3hqekYAeaejtd8fTsKEvtDXLM471BmlbqaXtLtb/EQFRJDsjLCkBYM5ZkHLKzCwiknIvihtc7saebOOY4BrRDQBIHtsQgOIPs64btRFmIEJ3xbDKhm30cpzzG9N9HLmSJlBF/jCelGtjt3HYlYAe7Z43hhy3hq5sb3V2V82+eFFGL1dVTgoizJr4xYdv/IPf/40vvnHjztHuziw2kXMezs7OhiHdvffm/QcPLPL7//wvn370aGd374tf/drO21+Qq6vjDz44OTkOkbdPIqzp2Z8/JvolZnXCq/CJ4/KZB208BZu/VK9yAL83Ifg1Uq8rNX8ErR8ko4VReRqhy/wBCdBEBUwBUEdDqu1O28tsM25v8akO8qcYipjwmWEAoCKr1SrEyMw787lnLiExIDJRIPI6xjU7CwDBzZ11DG8DBg5+064BPXDdgNctcGbZjM0z4eq+3fTKbcPUim65BH0BYJwiCACoYGeL5fffezRnm9HRLlnL/vU1IkWPlSMqIxiWVDYjtFD8vsAvCTPR3PWZBgzM/pjtuou2bZoQY2gCN4Qsklltv92/vT+/XF0OiG8dn9k0ZSdMmDDhtcREQE+YMGHC64U7bf9hf/sbe48iYR4WMKwAjbxumCkxhTY4b4uATdO2zYxiRA5GbDmbmiKoJEl5sVgOKWUVA8w5D0MyNUKKHIggBJ7vzNumYc3zwxv5xdP33n90tVhUiWxJc0c0QjSwJsYbN492d3cN6fT84mqxEjXRbGIgoqqmYjkzEiEYWRbJIm5QwIGlc21LWU5r8WQg95bIOauoZNGcR5sOP2qrZQyJaBiG5XI59L2XSPspDLcTZVX07ALMbfOATf55i9a5bmsBADC6417TIlb+YPy/Lo/qD9ysP7jJH40E5saeYWSPtTSM24utqj7e6PqGONhGwV09H2MXx22LbQhUqtLqp7cE3zY6PWz03D9ZB3HjSNYvE2jfrVZX56cnT242N+ez+cHNO6s+XZ2/6C8Xly/O6GbY3T148PCdp48fnZ1eINAX3vnSW2/evhyef/WN3ReXh8fPT5cDJKmC8jWFuR4gJDIp86TYN2/bKxSF8sv0i9nLr22M5chkrze6zvKsN71Gp26/jS/v3LSKf8FAEIXQnZ5zStc3xnUT6/X2y9dFFYHXLo2yy5FDtyJihhrTgGvHsxWG2eztxv/jXN3owrVL4RqPjVvnbs3lXyPxN0a3xDdsI+awGS0wfPPuzV//5W/89q98/cZus3940AQeVldnp8enz08ODg9v3Xuj2Zk9+8F3z55+tLe3f/v+W7tv3Md+9eT9H16ens5ms7t33yD6FwDXRNC/APiFOZDPDdcY5E+LzRDNdgsGJdOkxAy3HyD1jlKm9fUwSAkE1dYRoRSbRTADNYVaBXT8hP0Yz8j1Tj/mmK71ZZpOnzN8ZmDOslgsZrPZ7t7e/t4eIi5XKyCuOSvgJvlrhfL4ef9eZYZIbdMiko1mGGZu7G+mXm7ZeW2DQmQDlNoVJT8GMZsSERBD1QFsTR0ENbha9e897u8czg9nDC1ZAIiI0ARkIi80iEy2UVOAEbykRom0qOacwVTAXI6tKjlL13WhjU0Tm8ANAasZIDG3e81sNxha+KP/7p/8n7/1y/BP/9/P6+xMmDBhwoRPi4mAnjBhwoTXC23Iv9T2Fto3bh0NV6e9rbzkC4UQQogxxDZQjMQMVqSzqKJZNPc5Danvu26FYCp5cbUYUk5qwAE4ADJQVKKssLN3MDs83D3YD4EMIUN4cv7u//q//19PnpyBAeJ67YoAiApqO/P5228/aNr27Pzi/UePHz1+drlMwDEDJElMBAYmEkNgoiENFDg0UXLOOQ/D0Lat13YDqMYQSABY80ILvVkXPxYCu3UAI4po33VIJDm/OD3tVqtPt7K2l9bJLyu5qvUEvLThtd9sm1NAsGvr/crlvdyJ0kzVtenGGyPTZxsc7kYTNgpRN9no8RXb5I3XRN9IF2/uZi1VWrOJiDBS2LBWYY8ENL6CI12rW7eHaOuU4LghrpmUuoHL5XPqVxenJxezHG7e2Nndv3P3zaDWr5YXz1+Ywq07d+/ce5izPnv60eJqsVxc3To6eLjMV71ervIP3m9+cLwciqgXVBV0K+vWAA3RLbcBwBQ34gzXOrqNV1LS2+/b+qR+YlObB72pJdt8pbLHbqDtbiLlXe+4X5A4ultc2yNeW/9vmDjXfalPvfXwb35w86WNLl07tEoY1zjCBl/lBzDub9uS5trU2R6Jujd7aU5tEtC15fLhbUm9bW13uD/7O19757d/5etv37u102BgNJVutbg4O22acOONu83O7vmLk9NHH8wC3nzz/tG9B2Lw4gfff/b4EbZ7ezduIB9vBYg+Zn78HGI9QX6WvXg9YG6b/2k23B6ujecHbs+Qj9tszKdA3LB7shrmQaixPdt6OFnduMRi6wdVy1NH1aAW7QUEVSn2HVvpEPUCvX7fMBi9fKBe7+vL79pTkl4allcc8oTPBZZzvry82tvbPzzko6MjJBrSAMRUizy7TZYzyFX7rFZLR/hUjCHWR3QhoInYawAQlWeNqohmroSwF0jwghaqAipKBEj+dLneSzMzSAJXHZxfdafn5xalDzCP1MTo9ZmbtmmaACE0MYbIhAyAZiUoCWBmEmLY3Zl5GeCcBgBDxCw559ylYdX1oITAjMSxCRBprzmaN5rkv/oP/+2vfO+Hn+eJmTBhwoQJnxITAT1hwoQJrxf2Y1K2Jjaz3b1IqW0AkZAZiZmQiYgJENRMskjKmrLkQdIgKWnOaei71bKJTIigGUEZoZk1oZlTM6Mww9AAhdnBwexgv5nNKbCIPn10/MMPjt97dLrsMhJ5piaNlJQZAOzuzt9++61m1i5Wq+Wq61MWVQXRcSFtlnN2GY6YmgIKukt1CCFLFhFirnJMBVCA4hs7unOoltTRYRicj1Zwcw+TlIZhGPpe8k9u8Oer7Q3t5Mvv43rLTQlm+Wnbdgg/ejGO17ey7R+ANja4wR1XpsIpxC0++BW9LxvYtUY2GLvtj9gWmVc/sWUasiYpt3pu1xvd2Aa3yMRrhK4fiHklo75bnb1IjHJwdOvw8BCGdPL08fLqSlV3duZxZ+fmnbtgcnH67PFHH927/+DO0V6f9Oxy+atfuf/i6r3+rMvuevoKx1R3RB0PdNPl4ZXc0xZx+tIx/UjYKxreCiVs0rvXG17PNZ8FBoZAHufwpH3UlybQxqHY1ou48Xuhhyv1Zdd6tb3hhobyWnClRkGKZnnc51bQA5wxu9709sTZQp0pW0bWW82ua6NtJSZcP4OIEBi/8oU3f+tbX/2Vr7+1v8Ozhq1fdN1qdXVBRG8+fNgc7J8/e3bygx8Q4L0HD/bv3AWAi6dP/vq739uZzw5v3nxu/fHJiah+zAx51RG81nhFvOJVr5eXPg0j+wuHH8nLb0Vjtn+xa5vB9hiO/LJv4H+6/Y0YMEOINGtbAxARRGQidikroSGEwJ70A4iRg6gAAIcQOIjI+flFStkAEFDEhmJG9Oo7l73c182b90sxxpcOZfzAxz8xJ/zNwmPIZGbD0A9Dn3MOTRMCmwGoKSgCljq6iO5V5OUlVHXMHPGUpZylBjdKAopHL5yzRqJipwYKm0+YjRoOkrMaILPJKwho56XdCVqAMMad3dkOW4vq3wARQFLqcu4RmYmJiZgDBw7sOXNMiMhMTROJDIBjYL+i1FREc1bJptlAgImZox/mLEZKijZ876sP4X/6/E7PhAkTJkz4lJgI6AkTJkx4zUCmGdqD3dA0De/CLLrQGRAtZxAxNck5DUMahr7rUz/k3OeUJCcAUJE09AazWRtDMycAYN49OGp39qiZh2bGoUFmnM2xbRTIgLPohx8+ff/9p6cXiQiR0IUy1UzWAAAJdnZ33nrrQWyas9OLrEYcYhvEEBA5EBGpCJpxCMzcMICLcZhijE3bLJdLyRJC8BpoOWenuWOMUJc2zkMxMyKmlBExhOA+sSGErutU1ZdGP42BfgV9sP3+NjeB1/41fOlDr+R7fOW2TQRjfXtTrbaxtr+2PRhs2X+sWb6RlCt9reLStUR3Yw9mdQk5tv0yW+hkRVmRGlgdhsoRbrlG+zhsUBWjxG/NR740MM7CcAzNfHd3p1kuTkC6YVjtH96e37zZrjoFtdw9/eCvL67Oj27e3j86BMtPH3/03b/67hv3H9zYnX3l/q2ltj98crZYpbNFUrAqqN88EjOz4vECAKYbosNyFNdT1keqc/0bbJ7Gl/DSFPpY/gdeyc2OA4YbJQGpRAMMiRBJEMDMtWHe6a091T9sozWAUc2+Pls4/rkpdoT1Gd1QSZdYx2gzgs6e4SbLv30suJZVX38PwTaSBV5yItmaRWXst6IJNgZgcIMMXP9jzj7TwV77L/3GN3/zl95+697e7Ts3cOiWly9enDxadcPbX/7G/MaN54/eP/7g3b5f3Xvzwe7DL3KW5x+8+/677xI1b33xK0ph9eKjfrl4iTD/kRzl64mX70Z/W0nmH4FXnt+tcOMm71w52zIXyUsBlsKeGGMkQlMtdzlE13uOt90mEhLmbE0D83nY3z8EsGFIHDiEEGNkDsxETLGNzLRYLgmxbWcpDYDYNm3btEMaPnz/w+Wyc7eqIelymVW1aF1VVVVURDR7xTc1r6hrnn+zeWPzo8HNB5VtHOjLI3Od5p7weaEkjeWc+77vum63iWAgImYCiMKcRUTEOWjCIoe3tW+RP/FxM+C8pqbVv+kRInrUEwlMak1jLm5pUOKQamBIBOoi6PH5A4CAXqAYQAyEiJv24OhgjyVqLl8qVHNOOeX6PRCIKDZN2zSBOMYQYwiBmKlQ6gAxRCQztBhaRAJDFdBskoWJEfCyz1qKV6swZoZvf/sfffvbf/b5n6cJEyZMmPAJmAjoCRMmTHiN8J3vfDvrMGtm+3s7iAhiNgySkqqZaeqHnJKI5DTknLPklHISIUI1UMMQYmzjbD8wM4fQtG1s2tjOwnxOTYMhoBhk0WGQYZVNui5RmBnG1YuzdLWMYNlQKzNaJaOGAG2Evd3m1q1bq0W/WPbI7XyX5hyBWFVzHpgZDOazmYgiQmz3zExUEJGZY4yB4zAkYprP5k0Tu65PKalqjJGIASznLFJ8ooloZ8cX5GF0H3z2/HkW+cnWvp8kc/vEt7YcNz6WxcFX/LqhlLay1Ee7zn2WTbd9Mzb9lWsLhVdck77XeEBnjzf3vEVNb4ibvWXclnHbmocYvQ42uzR20dbmxlsbbDLQ1wj8DeIaEZumPTg8uv3m4eWji65b0cUpMyOHW3dup9328vTZ2dkpXF02Mezv7R8d3TLDk+OnJydP9w9vPnjjRgrz3/zmF84uu2X3ovc6m7Cti/eu11gFrjn8jbft2tbjr69Q/30ydfcqGxf7xD+33tj8uNbJoWZgsj5l19P0X256K6ZxfZd4/c9tEtv/XdO/W0e00XCdUkZrwtm3eZmCX9PEW1LL9cSwa91cb1Cccjc3GEsn4rXICSHs7sTf/rVvfuvrD9958/BwLwLZYnn14vkzETm6dau9cXh2cnLy9DhlObp1+/bDt4bzi5Pj48X5+cHhwd0331ysVs9OT64uLvb39ugXk6W1rVM+ocDWswuwZgpgrfFqZoK2ziuhDUMKBCCAg932xo29G4eHs1nbxPiVr3x5f3fn6vKcTJtAB3s7t28c3Tg6KI7NanuH+7FtUhYiiJFns5mnFXAIFCM2DXowhokIEM3TfQjJrzcyIEQRWVxcSRITE9Fu1V0tlufnF8vFYkjDcrm8vLg8efbsxYuzF+eXp+fLq1XqB0gCySCNN0qvGuoVGwyBwCvKqaoXgMCXLtQ6YhM+fyACeplkMFutVheXl/PdHc8eyzkDYGgCIBERVxfljbyfzRwgGGfxyFBDmQ7V8VnVwBDNaGO+I5hnqI0u0SiiYkagLrkuXx484uiX1un51bMX7Ts39yEEYiRG2iDHAby2oYpKGlI3DAzQ9ejVDZnJIzpEFCMTIzPuzHdijMzESLFhnDVoMKT/n703W5LkyLLE7qKq5nusGRm5YUcVUFtXV28zwxHOCIUvFD7zQ8gvwBeQz/yF5m+QQiF7RDgy00tVV6EWAIncYvHdzUz13ssHNTP3iEygANSC7C4/QEaEu5upqZmqmbqee/TctJmu1qtYgqstGNvyiH29Zzn22GOPPV477B/Ne+yxxx6vEUbVZFpc3oNzTXF6teJ6Sals8vKppiiSkopIiiJJVAWAiIp+D4nNIPT6PvRcKMCMiFzR994zcwKLSSwJRLEYLdUiVZS6qhK5gZh/8unji+cXmXLszAw61QwiDoe9g8l4PBpPr1bT2VKBnA/kAhCpKhFkD0FzXiSZWVEUapokEpFj570HQ+8DIvZ6Pe+9GWRLaGYmYuc4xpgzDeZLwdx4XkvMsh7Jcy0z65yLvxG++o63qLyvQd+8ioi+9eq3sZM3bDBeqsjtvbp3d1MJ2i0O+lUH2mWyW/a5a3/sxH8tK5gPdLuyv+1cdg6yFdki+qIYHp74+v766onUVb2aEeJwfMjeh8FkZCRSrabXgfjg8Pj45I6aTmfXm80S2N0/nPz43TufPb24XqyfXK/lVUbemOt6i0e9ccludiN7xV+7O34pMfnNeuSrd2oa4LeYV3y9cl99pC/qnrfVoHb73S6c0MUbXlWr/DHu3Dov3UUdCf2yNfXNrotd37tNpPd74a0Hp//hr7//3XfunxyNg2PZrJ8/exrrNDo8HR0erKaXm+WsPxgcHBxMJpPglg3GVQAAIABJREFU+OnjzxbTaa8/PD0/I4bp7CoKDCeHB4eHjffQv0J82UPsX+s5fwV0MZEm/ZmZEeRInjEAIXgC71xRhJOjw4PxeDgYFIX3jtDs6GBwejI5OT7qFT12/PZbb46Hg81qDhId2rAXDkaD8ahnKjkYNpiMfFHoTiCGiLLvAbKjEEwFDIDQwPLSAxVJSZAZEEBE1UAVziYmZgKmEmOsqmq5WJZlKapluVktV1dXV1fT+XS+mi7r+TLO1/VyXc2W68vFclWW67JelzF1vKHtPhANbmYCfZVX1Z9wf/nWkGXLBgCxjpvNRlWdc4Neb1OVokqISAQ71mCUV861L7sBBTsCerd07PyOui8DN4fH1qyjobZVSRAo6wbaeHVeaAXNo1oMFpvyar5arus+emJgACJgREBiQmaHBGCgqswV1WW2Sm8zEYIZpmRmqY6CaERQVxq8c469I+c4JwuJSVKqzdCxZ0A0HS6HAOkP0Ap77LHHHnv8TtgT0HvssccerxEI3L35Ix1t1vP54uKJ17ogo5zfTw3bNEMAiMiEWHjver3J4YSdB6BiNHRFAehABAzBe02S6mq1XGTTQJRsjGuqtWoyZFBeldUvPv7VJ58+FjBV0Jey6xHhwWRydHQUQm+53lxez0TAjExBVQDNOdfMXpCJGMyIGAzIsniFmLkoCu+Nd1LleO+dc9l2MISQ+eiiKMyslUITM6eYRCTGGFOK2Sr6j67C6hZQty+aN76gGt+0djszxd0Dv2KzrSK10S61+93SVnem0QivIBFuFb9b4O52twSqtn1luyLVRgB7Q3G9rcPNY5jFFMu6NgyT4zOWejO/SGW50Usy5WLcHx0MRpPF1ZPZ9eUMyYd+fzg6vXsOTNPp9Wo5PTwO75wN//z988vFZlF+Pl/Hl5j138KRdG36VVrrt9ItN7Tgrxu+qHJfeFY3tMyIXYdraeibqvrttrefHACvDIDYzg20Xbv9ynUB276+ew+abUslgjtH47/4wbt/+f0333hwOhoPVWV5fb1ZrUeTw97wQMTmz58g8uHR8XByxAjzF59fPX3CvhhNJr3B8OLFEwMbnZxMvLL75F81ufaa9tBvFQigAEaAhAygokJt9M0jFoSFx/Gwd3py9Gc//P7777398P79k5PJcBAspdGgfzAZjccjJk4iRfCekUFTXaaq1FRJvUnVWmJNCM4xlsnEOe9yPHWzKRHRsVNVRHLOabvooVOlxhg3mw0xAYCpiSQDKHwBCpYsm0Z75uM+8nAYQsj8oKomtaSYICw36WK2ePr84pPHn//8419+/uzFsxfTx0/ny02Kqt1okwxkJ6bUXpxtPPql67bHHxXdE1gkxao2tV7ROz4+ni8XdYyEqAaiJqqZKabsp3E7Ntp8kbz5VnaLzuL4vOMuld1WQNsMymYqakhaRzMyU7Tt6igD6NIvrKo4W26mi3XPehYoe9VkpbVz5D2E4Lxz3pP3fqB9QstfGjMHLZJijHVdx1gnjaqyXK4JwTv2nryn7F2DyIgwDMEPD1jQVmVYSdyTHHvssccerx/2z+Y99thjj9cFf/+3f2tpWffisNcrClcXzpl5RkI2AzUAA0R2zITERM57IESmMOiDgcZa6zrGGlTrclPXtUKTYabclCJqSMH32HlgNADC4IthJW61Xj2dLi/mC4VsMNutmwdmBjNCPDo8Hg3H69XmydNnnz7+3ICRHCLnXIJIW2VNu05e1bJEG6h1tUSknGldVXPaJSJSVWiXi0I+4o5UxwwkRRUFgM1mIynpS9OpPzxuzsNeUoHe+Ah3/jXbvKSH3uqAdwrE3UJexQxv38PtVK/5/MZyadwSxa0Cus1P1Wl+b00tb6qErZtL3uAiG1rCtmbJLVW+TRzX9p0dsdUriHo1KDfV9fV0sVgNR2F8dMKk68W02mw02fgojI6Pil4gWc+m17PZTJGP79w9unNyCCCA8/lsMb8+6o3//L3z2UaeXa9/9ulF0q/QMb5e3sivt+0fpVt+o4N80U5beTv+lpDKzbyWALBt4m2X3tn/VsRh20leVSpAR15Yy2nf1GLjNuDyEnqFf+fR2X/4q++/fX9ycjzyzMvp/OrqcnJwcHxystmUzy+eQV0Oh6Ne0fe+t5rPPv35L2K5OTm5MxoOytVyU9Z379/Hg+PPy2fT62vT3z3H6b88bDvBnxIyE6ZqjOAQ1dShHRTwzhuP7p6dDvrhjQf3Ht6/ezAZDXqhF8LhwWgyHAz6PUfGaCAQvBa2xsVGkZgIa6doIinWZaqrVFemMWcDNrO6srRMCsbEapqS1HUtklQNAb0P/cFgtVpUVQmIrQ8uqWiM0Xnv2BGRxiSSBNA579gJoJipNoRj7bgZ9kHV0JDQhR66e2Me4vBs9OCDR0fLdblcVdP5er7cLFbrZy+unjy/fPzsYrpMq0pj5uObUFF3k9/qG39yXeXbhlluFgAAFIl1XVZl2R8M+v3+utyoagghJkUVv00F0Tg83ywKtwk+bry58wI7T/4u90Nzt3SjPhEicgJ8RUaOLmCIUEaYLtPT59O0cCOPReGzI3p/0CuCdz6F6ENwwTlGYDNEMzQ1RQQk9I4c+17hDHrZzDzGpKbYREZz7gR2HLigUPQG/SKAi1V9BdEY9zbQe+yxxx6vG/YE9B577LHH6wIbrXE50uOrftHzDoq+d0YOkYgBuZk2EDt2BMjEPvgkMUkSUVOxWFfrWiWRSVVt6qqMMRIhM0tOWM4+OHK9AorgyMxx6I/rRVrF1Yv55npVKoBlz4KGmcKGv0Q6Ojwaj8bL1Wo6m01nM18MmRWRVCQT0KoKgIjk2CFCTLWqQOPkioTofWB2ZhZjTCl573NKd5EEWdHNnD8lIudc5qZFREVADRBTXYskU30VlfXaoE3e9hKh0+nIXkUud5+8gqS7ucH2hb1yO7yxqWFDFH5JuTek3TvHuqU63a3AzarcMgjF2xu8EjHWy9lsfnX56OCsODopBsMwuPrs459ulrO6Aol2cnZaDEcHd+5s1ssUN5/8+uOEPDk8Pj3vofPPPv+Mke5Oxj957+7FdP3s4mq6kfi1klN+HSH969Thvqgu+NIGX4Uksu1vvPnH7kaZjMLbbzULrW/Qw68+6Csq/UV38as2/aJiEeDh+Z2f/OC9H3/wxt3jUWBdTK+vX1yqwNndcyZ7/vnzyyePD0bj/lHPhX613sweP15MF3dOT4+ODsDSerW5e/+NwdHhaj5dffrLZ48/6VR+f9y1FrdO8Fvoca94Dry++NpLDtqzuhE/REBGcMEdTYYnB5NerzcZFCdD/8H77zw8PxsO/KMH5w8f3Ds6nDhGSRFEQJNpkrqWWJtFjoCC2YUAiYEYwCRFTTGlGOuK0JiQMItGJaVKVZXy2CcaY6zrGKP3gQsxhLRaxXKDTFQE8EERwMADsJAzIGY0FTNVcYSeGcFU1VIiIjIyS6Y5o5wiEhIhpuCC7xUDDqcjJj5SQBGr6rjelIvl5vGzi0+fvPjl4+cvruvrRb2o6vlqtViu12VVJ0mK3Yi7MxT89if8Hr9vbMdxVU0pVlXZ6/ezjbiqWoNt/NrMcoq/l8q5Oay3Gzfk8naU39pGN2miVaEtERG5iy+/6iAGoAi1wKqS2bLsYy+gN1QEA1ADiCkRmgsueFcEH5g8gid0TMzEjAyMjM4xEyGhgSloEhHNiUHMVE2VyBN5Zi4cB5RR6AWCguzzQygWv5eE1Xvssccee/zesCeg99hjjz1eF6ATvXehJYJzAPWg10dLBMbkvfPOB3QOkcBAqlpSqqtyuVpsNitCZAICWK+WmqJjIgJVKcuNc64oiqLXcz6wK/r9oR+OcTwGz+Y9huE8Xi+rz2ertCqlE9h0JKqqmAE7Pjw+Go1Hi8WijhGJkAkJCRAYARrfZjPIbhtIKJoADVu3ClPNTpc5YY6IjEYjIooxqgoi9vt9772qXl9fE1H3sq5rTaIi2ZTDNKeVe334wFfxbt2Mbmcit72yYDlLz5cVZreZr4ZuacSgneHxdubX+S7aLWqmmWzeVqa2/Li94oN8+M4OoUkud5OMbjXXBl+kmm1mqdZq23G7S66oqcTNarZeBB6PyYX+6OD07HxxdR2rcjm97PeLwdH44PgYGaeXV1W5iWWZYu2K4uDoTrmpNvPrYPjosP9vv/fws+dXf/fTz69X1Z/wdPOVRMOXk0QvkRDwaln/9k+DL3q1C8y9BbvO2ZZs7QFuKqot6+qg8RfqPsedmwi3ZPc2d+a473/84Vt//aP3zg56AXR9dTW7ulaxew8fONAXT57Mry8D0+FkMhyOKNZXLy6ePn3me8OT+49iLNN6NRiOBwcTq6vrZ0+mly+Kwt+8BH8Elu1leWlzyn/4Q78Gh/wmwFsPrK+8g3UdKr9DJgW540nvBx++85d/9sP333nzzft3758dj/qhcGhSpbpUqV1cxFW1Wi/RDCRJrE2zynnjCL13zjkAVDFEAjDR5JABTGNNjpm9mYIpoQXnEME7BwCqGutYOa6jGwyGIRRM7PlAbYxEoQjeubKqiMiHYGKiKqLc6zExgAEitauIckyXiFVVNOU1Q0SIjKICkNgAUT2boTp2XHgbMBwMDOl7771RCixruFpUL66Xj59e/OznH//Tz37x6eNnV/PNWk0aTXTzsx177Iu77h5/UGSiWOuqVtOiKER0vcmL3lDtC75dwK6a+QbHDC8tHjJrm3pXKa0qdQ05PkeUzS9M1bD7TrbzBaTtKgoggAl5cHB0dnKY4kZTrRIl1bEuVRMyMFPwLjAVzEVw/SL0e70QPBGpKFNOC4o5N6jvFYaQ83LnWAuImQIAqkqsS8UeqcakB59TNfi9XfQ99thjjz1+L9gT0HvssccerwssiDPmvu+Pxj2ooXAgEVWzoWOsSqtMUoxlralWEQOsqzLVFWStMoKKIgIyk3PM7AYTH0Lo9cOgz6FA5xwX5DwSSxVlU6G33/z84//r//y/Ly6uVAFb5siw5aANnKNRPxwdjIvCv7i4irFiJsyboIIpETrHIgI5QU2TUYnQoEuqbmQAjUjHucb6OStY2BEhGWhKUVW9d84xgMVYiaiImEpMsSyrmKKBfk3p28vT42+samzZ9O1L7ObjdmODHaOHG14WmX1G+xIO+sbp3RIpt8zdDe7lhsy6/WzHIuPGyXYVe+mjL+EqbafMhuXuqmQdT90lhtw1ZgDEXVvg3SMSAaHFzWJ2oVpv+uODotc7vHOfKMwuXlSb9ezqogYZHownh6equC7rq4unq9X8+Oz84Oj08OhOvV6Z1EPv3j8b/Hd/8d1nV+vy8eWqbgT1AF9+hW+e01dAl5Bz9+XLx8KdGfuXuMW8XM43wFco5Baz/HKYxG4UBNttDHc7ITbPhd1G7N56KS3ly9R0J5K23auOL22ze2ptpKI5xd0gigEAEMB333nwF997+/2HpwNn5XI5X67Jh6OTg/5oMPv8s+sXz0DS8cnR4fldx+7qxbPnT18IwKO33+/1BptFZBf6w76upk8ff3Z1PeWif3TnjOhTgFsuHL8LMftb+9frQOF9u8zzVwqT4I2W336EO10ZkQDITLp+mz9p6OY2v9nBpHd2fPDg/Oz0cHJyOLl7cvjo3tnD+3ePD0ajnvOyhJISqsRKpDZNq5rMlFTAzDSZ1ITInjz3EYwIgncAlBWZYOYgBOeYSDSoGoARcs41KKqI4H0QkSSJfCjGI2ImIAQws4AFIiA1NrjkPUIeVQkARBo5MiERM2arXFUVJe+QyLISto0wIpq2F0JFVbXh8QBUDMCQoHA8AB4rHo+K+0eDN+8M37938Fffe/vyev75s8tPHj/77MnT55fT+SqVYpVC6m6PZkTqFLFtq/yWZ9rr0OG/HF/ldviq48bvVJFXPSNziapWVmWKkZmLInjvJSVDBEDm/J3Rdr2esys0vNQ6CNYG9wDalJgieWjPX18QEUVFDQwJmRBzeg5i5kSoiIa4jZrblohGAAXYRHlyubp3qtTr9QOikCVkcwhqlr84GiCgmZrWsVZNdV0RsXPOO5cP5Jzz7Ng7H5SdI0fMgTwhosSUYjKDlFIVkwpHlTql6Dzq6KOPPvroo49+x1bYY4899tjj94U9Ab3HHnvs8bqADCWG8WEoej2voJAAwCyhpVhX1WYjKca6rNcblQhmxJQXISIiEAJxCIF9cCGQCxwKV/R8KFwI1CvQOSMCBU1iVVmvVqmK4Kpf/+wX/+//83dXV9NMXqI1FDRAY98QPB+M+5PJ0Dmaza9VpegFIkdEAAiizByCVzVVZc7TBTQLmWxtEqY3izuNiJzzRJRSNNOsBUNEAEspmllRBOZMQMdsD22mKcX1ehVj3VCs35x9zmbT32RvBIStHKid17UzN+u2aexqm8l/w1CbQuNssjW2aHxvb7Cat476RVPcncyCLYH4BfXf0ZluM8ZlGNzgaLasddYZ3VjK21pCbnfuLuLNMnY/ak82/wZs9XMGQATOu6JwZLK4vtB6baZFuOv7o9ERSIyLq4v57GpZl8Q8Pjw6PHXrsppePFstpsw87I+Hg9HxyelmOZe6GrP+5N3z//rxvatlWV3Ok7aW4q/Kv3TjBb7iwn0Re/Kqbb9ws46tfmVp28CM2Rdt88oCd96E3XP5SnV7OYDSaNLxZmnb+MZ2ob21OvimQduOu7vHF0WG2h1yBfIPvJVu8Hbn7IrCxs8Wtt7vmdpwRONB+Dc//vAH7z04Hjgp1+vVQl0xOTkdTMab6+uLZ09jXY8mk+O7d4tBsbyaXl5dJJOT8/O79x+url44Dr7ogabLX//q+fOnODo+uHNvOFki4cv1+Kb4KrfzHvAl4a+XtsEbPb+Jlm4HBkJSkHbVRVOIIyoc94Lr94phv39+NnznjXs/+uD9R+dn9+8cnx4e9INjMk11XS7W81VyRGgqkRmJUUwcuxA8AIiZkTp2zjnnWFVUxTufB0QRNTPKKXaZzbSu67qucyIE51xSAUDnPYqAkAE4731RSBVTSqrKjpgQDNRUzdg5MzDTzGCzs1hHFQEiQAQkAAAkJFADU818oiG18U5AZoCGulYzQlAVFZWkmVzkxIgICgP2g4E7DP03T8dKb9dRnzx78c8//+U//eznv/zk6bOrzdU6zco4q6p1FeskBtC5cyA0SZJzZtEvvmde/7vgK7LPX+VEfg/s8ytGqPzTrNyUVV0DQghFEcJaBACIkJnyM7MloG/ERF8eE1v/NDQz53KaaAPDbJIGeY1bAlNjFxqNAWd5PQiREaoh3FqZ1n4xMYMyyvPp6npVlqrjwIV5StJ37AgBTNASmIFJSpKSqZhqTNEsUR3zWgEE9OxD8EUIKbAPzgUPTRZCNkQiMoMoUsU62hqI1QDN1sfvwfPnv2Mr7LHHHnvs8XvEnoDeY4899ngt8Pd/+7dQL11RMrhqOa+rRbWcp7oCEc8U66rarMEEwciTAlpWLBMSuxCKotcr+n1fFBwK8AU6j+wQCQ1ANW42IqIqlpLFlOqYYooJE8bLi+vLi+uyimq3ScZMrRZFcXh42O/3AXG1XvkQTo6P2RUiklJSMyby3vf7A1UTUSJm4sGgY4ssWznnmU/2ekbEuuZsEs3ZMQRAkqiqa/hoyDQQIWX/jRhjduHIZO43nsfu8BK7efsAbq02zZxYx8zlmVzmYREblhapeze/zrshoSFhs7URGJi2iu8sTmuSQ3asdLtvKx9uaDq4bXDRVSd7FTTs4S6BeEvx+iX0a2YPoE021W5h2NSnzWvYHqAjG7ElGHbY7Z3iOyfJ9sOWBwEF0FxxNhv0++PxZDgapNXTzWoeCl/3e0IhFGFydKJJLi6exvmVLwIQD8aTew8eQapVUr1aPf7Nr+8/evjgwaOry2cXT5/E5XzU93/zvbeeXq+v5utVlJ1r+AW8OQAAaFYHvooleFnI3EVTXt7sS3jkrnluobsdvkRAfav8nXd2JYetwK3Vw++c93bLzCYTcddIeHPr3FtbDbs1N0fbp0y3Ld7qoq1jmmzHMgYJb9QB2/+a2gEAba/JTh8G6DJldv8MAbS5d0RFd9mTQc9/5+17f/Pj77517xilmi4XVbV58MHD3sF4M19cfvLrslyPJwcn9+8NxqP182ePP3tMYfDorTeOT+/W08V6vRr2HGmaPnn+q199fHR+Pn7zndVl2qz/603T1G9XGvxHw9cI6/0RYbu1ah8m+PJH3ecIhia55yAAt8s3Dvr+7Hj0xsPzD957+3sfvF84OxoPHp7fGReux0iysU1Kkkwjmw69egZmQCN2RERqnDWYgCAOEzdVAVM0zVYayMzsQuHBIMbaJCZNZqqSTFNZlUTkgxdRAIjMRVH0vK/rul6vNot5zr9pAAmbmCsgEKKqAjZ+V3nQSSmpKFEjuGZmU0spRRU1Q8KUHavMMk9IjvL9VW3KFCMSMjExERIAaH4KgaEaMSNQEnOhH3oDYH8y8j/5/jsfvvtwsYnXq/qT59cfP37+jx//6tefPn/y9DqapZ1BgG13uctO82zH2a/I2+7x26Gq681mvV7HOjrnfAi22dhL1xdvBY/bASW3jnPOzOq6zrRyfhbnLyoAgACNDJ8QwDPx7lDYrlFhQAbK3mhtOL4LT2cnaIAIcL1eP72+pklwHjyCmZoCIRTeD4oQipBLzLbOpgLaLLBKMUlKkkQllZtYVQagBkacXUCK4H0oiqLfD4Vnxxr6mMhXVQ0K//APdGf4B2+MPfbYY489vjL2BPQee+yxx2uBVGzcbASnVwEsLq7iepaqDYigqTFLSgoKYERMwfd6PUSwnOOeXH8wKHr90OsxESIaoohK3EiMJklTqus6c1iSoqSUkrHvAYblqryera5nm6xmwhvkVDMDGQ0Gd8/vsnPrzWY6m1eliLJBtEw2ialajAmzFCtnMYSckxCgnatwFmEBAAAzE2Vljcv50PP02LHr/gYA733+I9Y1Ima3aLCsuPr6k9hMpzXWtAgdlby7ScPJAREh7VBzAERIW2+RPCMj3OFmibJuGBARCQFzCZjZZ9CWRNtqwfMPa7hrIsItEd2RLFsqd/cssg90XlDeVhpfItWbaSbunhvsME0tBd6xnx1haK2EG6C5Gkhbx+d2T+gsKW5S35mV3GFjqaGvTQHEUAHARA4Oj45Ozk7Oj2xqWs7KxdWTzWJ8eLd3cj6ZnHjqicL1/ElVTmdTFEjj8eG9B29dXLx4/vRp9eyJxtVb739nOD6oqqosn2yWlx88fHj54++URv/46+fsPTHtVOvGVdlp9yZHExHlC5P77dbUHAAQDUy3BunNBD5vk7fPHSKftZoiIBNpox27zbk00/ud4AdmQ/W2dGsKJLWmyyAAEpq176vkvRqZpKqamjZ0dkMj7DQINZESQOSGKDfd0t87wRXr2g8ghw3y3WKA2xxVLenc9jCwNnjTdrCmx7V3R+bMd5Tx246ee8+WfW67YttSZkkkpVjXdazrlGKuoWe4ezT8H/7bv/zgrXsnh6PN/OJiOnvrjTf8cDi7fDF9/LnGdHJy9/DstNfvx+Vyfn2xnl0fnvWL4GIsXzz5zbBfpHL57OLp8xcvzt987+w7HyQKm1/9/Or6SvV3MRL/okfTnnf7crx0nzYUc/f+9qPmCQU7zZStl5u91AEQAAM8un/n4b0752end45Gd46G986OHt2/+8b9uybRMw4K78HYxCyZJSMBVDAFUwRBMUS1mJWdJkjADAiqppKg7a75BhTLowsWvR4AVFWVddChCCoqdVWVFQAk76FJESgbdkyU47giQsT5Wdqok1PM9LGoEiGzy3kOmb1IUlVCykSz8wEARCSJKBgSaXuPNsMRc77NTA1VJYrmXMHOGZiIdHSiKRExk0NIkjYgNbEfDfx41DtBuqd4/uD0zbfOv/Pe/c+fXjx5evX8cvrs8vrZ5fVsUW/K1PCCu4QzbIOm0MRuX8M4x78U3Aj2mkFKsSqrzWbjnev3+ovFwgCIKedzbr+9vLTkq3se51HMjNsvNZS99VXzSOLYtQ9qQ2zcOfKOqiqqpmYAxGymhp2Nx41oVr5Ra4Dr1frJ5dXYHxZGaNEIjckzsRqqQVJ2zjlCcIRI7digKiZi0sbvQcWiaBIRMVVNsRIQZ1Knek3kiFnVDHssiQGK0zVW8Q/bLHvssccee3wd7AnoPfbYY4/XAyTl5Hpo2ne4uJ5WqxmBOUZiNBB2iBzUkJjZh/5w4JyPooZMzvf7QxcKcE7ryupKY12v1/VmGTdLlagisY7ELvSKKJLUFNxoMAY3WF1dzxblfFknRQC6YW9hzQRgPBrdv3/fDGbzxXQ6r2oTY0D2PjjnUkqSdVfUkErOOSKJMebpTdY75/cRsZNCNzNdx3ndMQB4n605EgAAomM2s6x6FpGUokr6htPXhqSlhsggRCQkhlaxk9kyaoU9zrtMX1KjYwZmduzy6TATs6OGk21049Qw0juMdUMqG6ioilmTNSdf3E5P2hD0xK3nZ6sNbSWmLQvd1rMlrM2wNTXtzqDj9aydYGYuGVu+HbdFdYTiTns3FLiYaQ4kNNPSLIJqC1VTM21kucTUlNwyjI1OVVv6ErtLpWaioAYmdX14eDgajYvBmPRonVZltcQUF7PLfjGEPrEPd+8/MFfN51eL2ZUZOqTh8PD45ExiunqRZrOrixfPRgcHw9EQzu+F2XJebT5843it390IJw7Od5PnLa9/u0sAiAiA5c6Zp/QIyI5bcr6x0YgpqoiZETMAqIj3ARHrus6hCSaynFUsRkQMPjQJPJluHb2O0cxySMbMVJQdBx+6DaxxqnEppWxEQ4jE1C0gSEnMlInNNEmKMaYkqoJIzNSx5x11l9/EVsZuYFll1jZ4F8PAVppvrdIttx/nm6OV8FtWjiOgtVxgF67JWunscp4jME2vUzXTHZdwBEAiyn6+ls1zdYejbt+NMVZVtd6s89MATQEWhhIiAAAgAElEQVTtaDz84bsP/92PvnP/7ECtqiQNxpPR2Vk5m149/mw5nY5HB4f37/d6YT2fzV48q6r6/N75+PSMQNdXz/seHabnL57MF/Ojs/O7b7/X74+eP7+cX7yQVMMNpudrSYP37PM3ww1mrX0n2750Clts/zcAvbXgP/dibjtt37kec5/5b77/zr/96x/+xY++f3YymQxCzwODgMQUKdV1XS3JjAAYDciQgIA0r7ZJUVUM8vIbaQ/R9FUzJUAzUG3MkFUtxSgx9vt9RKzqWkWYeXJwYKqpquJmo2biHIKppqquYqxVhZkRCQy5eQRZSjEvBmJmZjaA/DSIdQQAHwoVNTVAEBVR1dDDhhZUADBEZibH2T/BVKmRoVq/12PmqiwNkIhDVr+qMTNlD2okdq43GIhanUSkBkuGCc2RD6NBbzw5fPPNs7/hD8uqns0WP/3nj//hp7/4L//48998Nn92uVklqURqkd3GtG3DdQHQPQf9DfCy5B9MLcZ6tV6PRqNev+ecU1MkYuYuMppH6ls75sSV7RjX6APyYJ8DtDnYnr+8mWlKkm06mFlNJYmopCSSknfMzKoJNDtBv6JxswJ6ul4/v8L7B/0BsGqVmHqOsQhQJxWLWIfgil7w7Mg5753P+gRjJmTqJPtWSRUlqWlV1VVZlZsKTKROm0XFzEWvF7GMYew1CdPQ9eJtQ/899thjjz2+TewJ6D322GOP1wIWojcAdqoWmP2g773LBKL3ARDVgIseuYDEjICA3qyOUqd0fXUVU4pRQCJoQhVUQRGUmNcjM3t2jikMhj3yQcCFg9O1+Onq2XRdlYbIngFFpJvjIAAaEMJwMDg7PV2vNy9eXM4XKzUmCsRYWVVVlUimvVxZ1qqKSM4xEUk7C830k6qGEIioqqpM4xJRw79J49eZibOqqpDIO+e8V5Gqqkx1vV5D61F4Sw33pcDbfyMCEnKezjC2MmaiplJ54uV9IKaGWAPI2p9m0XKzSU7Eg2atQBVbQw7KfMKOALQ9WdiSe1vNcXv0RnVN2dlzx3sjy4lhKwVszaiNOgIaOytf3FJ3twhobGnorao6M93QvMbuQqmBttLsHV7eMrncGolANonMF6VlzXdPEjpac7vsV8w0ywmD9+wcMxf9oY4mIrGuqliWi+mVJOiPJ/3R+DDdLes61lW9WU0vzZR6/eHpnbuEeH314vmTxymWRyenh6enCbi8nJ0OwnfuHTx/+8HPnlwrOx+KXQGyWUM373aREAoEyInCADJxrCml4AvnGADqGCWlIvRu9a2iCPkqOudDCJk5ijENJkNiMs0m5ua3PHiDXm9ws/9i18Rdg+frFkLRK3rQXls1RUTnXIxRRZ1zBqbaKCg77TZzR5MZ7PDI+UAGRl0cYqdLbWMX2+4JmHOdERG5HGPIOjRR3emKDVHfdNeWgO76aRNM6UIXbYfLHX+XgLamFfKtomZmiGzGIl0cCwAGhX/v0d1/9+PvvnN+WDiqIw4Gw95kJFW1vLgslyvvw+HJSa/fq5azxdXFcrEgdEfnj0LRK5erejZzWq/WVZ1kcHzn3lvvDiaH69lsdfVCq3Xh3NdhnG+h23HPOP8uuMk+d8DOLijLe3d2yJpNsINh7+x49J133vjw3be+9+47988mZyfjk8OBg9JW8woSSLIUU11nkldTAhUzSLFKqS6CR7AUa5FopsQkKYmIbRd5NFxqvokyy8yOVTTleFGMeSAzs5TSdDqVlHJQipnNtKo3KcWsH0UkosbOAy3nFUTPzoKpal59kt2lEbEmBsRe0W9uFgRmdt4ZkKmJKQAaWmOpQdykbyPKi4cQ0HuPAIzI7LwPzE5E61gXvYKdUwAxA0TnvENw3tQAmV0IqorEvmCxlGKEtBkSD4/6Bz98/ztvPvj3f/XnTy9Wnzy5+udfffLPv/z1rz99stpoLaAAaiBgW6X6q8yI9vimaL4RSUqEyEiqWlW1mhJz/mqFTVfEW7tlhlqS1FThjq7ZAHKfSSKmqaqjY2dgKaUc/sxrVFpTtbZhEZDIiBv1exvhhvZXHnQrtTKr9IEMqIopxWpTrR07x+yIQ/BVFRw75zh455i848I77x14RFNQMBPN5hvIoSgODg4JUUU0JWvXClTGJfZ6E/hsul7Vyo7+1//5f/pf/rf/44/YNHvssccee3wh9gT0Hnvssce3j//0n/53WKAlKHpjXzDDGK3nnVdNphacy7wesDNAVYmx0WNWdazqvDy9TnUyUARgRkfs2bH32TvCucAucAi94cD5QgxpcDSfVb/69OnTF1fJwGV6sVsy23BPWHgejfqHB5PHT5/NFysRcN77UBA5A1DTnHmpyYlO1Ok6W2aS83rh7B4AjeAUWvsCE5FW+ZtlzmJmppJl0Nn6OdZ1WVamujP/h69G8dyiqhEQgbJlIQMRcpbwErfa5kb541xWL0NHs2ZxEAI0iQXzdL+lh80QEA0J0MzQAAwNs58yIAJ17LBmFrelZtuSMdtcEGTra2vJvewQ3ehWb51arl5L8zXsMuzY8UKrmG655I6E74iATCtvNWlmjUEFIdqWswZoldjdIluEzMLsYussspV4Y5OCzgDQEMgMDUEpmVqq61hXQ+dHBydIbjm9tqqcz65FAR0iw2ByfCxSLmf1ejW9uKwqPTt/MBiMT8+8qV28eDxnKHq9UTEoBoNJjLSx8yF9/9HJ08vZrDGVYWwSKgIioDYkaD4xMyPI7LmoGYARcqfa0zxvNwQkIjZrWCFsLFkZwYg9s0NiUEViYiBmRFITzFRwjkg0F8cAgNkhoWmzWp3aZfjdNQQwMdMojhmd6zhxbHxhEGFrAEOIZNBoM8EIKWulrbFKbxsVIEuYsTUPgdZ+BJrsYe3Rs6y/7Sy0Gx8ByCuvsx8IGAA1qkZraWYg7HJrtnpr6PqObUMr2HY7a2rSbtLS1a2zSPcZAgAw4YO7x3/xg/f+6gfvDZyKpNAbDAc9F9eL589Wy2XwxeTw6OjOWb1czJ89LZdzh+QHEz+YWF1pWcb1cja7VMTB8Z3Dh29Mzs7jcnH15LN6uSo89wqP2N5af1r4WlrvPxxs5/9b72cO2hCNWqYrP+L7BR+M+g/Pz95+cOedh3fefXTvnUf33n14D7VCrWF9uSnXdbkiMJOkdW2qpoCAqqIiahpjnVKMRUAETaKaAK27lQyptYgBQCRiark/B2B5cQAAOS/tCoacJFDMFBCdy/FXACPnGTGzzjme1BgqIRMxt/G8zAciQl5tAwDEHpF6vX6OJCWVEEJRFGJQx1hVlQuemVuXKWTnnGMiTinmlTfMjAA+9JrhjlwSoZp9EYjZCPPyJCIGRHaQRJAoOBIxQGMTk0Q55EyOne+NisNh/+HZ6WITX1zP33t0/N7Do1/+5uziury4Xlxczy7nm1WVIlirV2/iYXsN9DfAK6+ZiMa6RsDM4UZE6wz8kdpfTUQk/8zPNUIEZgAgpCydzgx01t0DooqaQV4KlhM/ICIT5+ggM+U9mMBMASypylb8vo3Y5GorQC1aJjN0xJ5Q2+eNqmgUjRCrGKmscrpO79g7Ds4VwTvP3rFjQgRDI4fkyDEHdj6E4ByYmgphk14gKBXc61F/Wqd1LCUMWX4XV6U99thjjz1+n9gT0Hvsscce3z6KVarGzi/CcDTpjwOMBmAJDUETiICqSdJUl6t1VW7qsqzrKsWomlQEVB1zQPQAQIjOuVD40HdF3/f75AJzCMWAQwE+IDEAOlHgwWrz9P/7Lz/91W8+M7NoAgAKiq32GQCYcTQsDiaD4bBfx1hWKRSDwWjU6w939WcpSV3HwWDgnGPmuq5jjABYFEUIYb1ei6T8MtM63vsQPLRmuEXRyyrR1WpZVXUILvNxxKSqzrvryyrWlarsrCT9aiLoxnPj5jtIgGAIhqDWsLGGZIBqhmpqIBKRkJh2BaSd5XPL/wEAUKs5xo7Dy3xzy/EiICFya66R2YwsIN0lEM1AG8Ja8pXZcsRN1fPEsWPpAAA7n4MtAd14djTqVwMAbPLX5TRWuyVulbmtFDrzfmhwg3227SGze3BzYhnaBhA6AW1HPOIO7bgV3AIgithmvb6+upgd1wfHg15v6FzhXbGcvri6uEimAmm1WZ0/ePTgwVub5fTZ40+ev7jaRCkGQx96/cHw0VvvEEpVrS9fXMzX9f37j/o+hNnKLMY79Muz0d9/vlit1z4UiCQqmehvnLi1ccAQURLBVqRvZkmyMQWVdQSroWXZxayu67quvXOZYo6iRIjESS1Vde7bxG69qW5YyogSQWaZc4OIWkcwmVl2d00ptjYglunmLKUM3gORJCnLjWuW1deZOGZHmcRNkqzNFqWQJ+NiZq0pDqTURH1yr9BMB7Wat6yJ7u4T23GGQSQDVTUyy8RYVkB3CTVBOw9nUM2y5ZZdwq7lVVVvqP9bUT4A7VSklclnrxqR9kCaUhJtzqgX6C9+9J3/5i+///DOQb1Z94+Ph0dHcbO4/PwTLUsVPDw5Obl7JkjPH38W10vHNJkcHJyey3pFUkMql/PrX/zzz9773g9P7z8and6rq/jiN7+5ev7C9wf9/iCzNrjDl/0p4VvnoF91dIOdFJYGoJQfmwgmhgYO4GwcPnzv7v/43/+Hv/zRh9996z7GMq7m6+nj6fXFZj0HtLqqUl2HIoCK1NGzc8T5kWjQOGkQoqaY10nknAWi6pxjDoAMgGYokgDJew+EoqpVhc6h9yjimH023slpA4mYOKfYJeYiBBFZrdeD/qC5s0yhdaaC5jmdnyhMHQetmnLIFgl9IqSi3yNiVati7bx3RUGAEdblcjPqez/oO+8NAPJ4AgAARdFDRFBrsxhwSklTZHaoakxiKmYOGcnQMmNJBqBSgYC0i2ZiTADGgIgmMdbrpaghOeeKsfPj8/E7977/73/ywXy1+ezz53//01/83X/+h//8T08+e7EEgAgmeV1EOw4CwJ9ejOeb4+WATB6NJaVqUwKY974IAREVjJnzczX7MhG59sGrTdAxB94p+4wRMe/GKbN5S/6CAbvfE7YHzj1Cs1xAUqxqsiRicYd6vslBIySxKhq6wKHHCoGCJ3NomlKq46aqYh3FwLLwn10WQaNBXn3mHTERO+oP+kUv+GA9oZQgusiMzOSJDAFRkTA4Gk4mk+vlxaLkOtW0J6D32GOPPV4X7AnoPfbYY49vHyn5g+dlHI+KojCVVG1itYlVlJQ0RVMBVVCNdSUpqgkaOufBWKA2TP0QnHfEDETkve/3KQyo16feEMkhEKNHIKgTSFVV1WK+jlR8/umzFxcXq/UaAEwkW/Zaq2hEAGY+mIyHwwEgllUUgfHkUAGqqr45GUJu58wtrwQAmTwSIgTgvNDYzLz33jtmzpJPZpe1z2bmffDeI0JVV9myAwAc8zVYSt/U/XnnlDpiLctu1AwBDEmTEsmWb92lkrPrriNsDZJbpXIzJaPMAbd5CbdO0s2FaX60KX4a0ZA0a1dzmdQBG7dc05xrEaHzOchn0gppofGHth3iu9katrLsTu/czCE7PWpHjrdzy+ZcIdOT+a/uo85BoatFfr9tb+ok1bunjZ1e0CC7MrTpqRARNVaiQVO1mD5f8rB3cjYcjBw7M5nO5kljuVmkFNeLCdqh98Pjs4cJ/HIx3awW184fHZ2ORqM79x9dPn8yn12n+nLV64+Ozor+wC2nQRY/ePvOZ1eLq+eL5XKNRE2yx5aDzguK872SKU5oKVdVRURmFpGG52XK9HFed1zd6Odo26Zsmj3GaJYLcUSYPWqIMC/D78w3cwWwMVaGLHU00xhTkyawcXym5WopIrGuQ1EgYkox25EbbNslpzFU0yypzhbdW66ndVzZSXNpuafd6g/bTout/3n+kbt5TrSYY0HWNug2QtJUZ0suYUNRWOM32lbX2g6ZPaOb1Jz5wGZ5bYWqaJNfMYmkmEzVOfre+4/+6gfvvvPwhJyRK3rjsSOIMRpSpXB67/748MgAls+ez65n/Z4fn5yOJwe2WWm9Ltezq8vn0/l0cv7m3Q9+PDi/V1aby9/8+vFnnw8Gg9HR2Qjr8fiwvVm+MRX7L51Wex3U321CMwTMtrRmuI2PGgKw4ZtvnL396N67jx68df/44dnB2cHQVhe//qenXpPWZb1ZqERGcOzJcTLnmJHIkIIPPiuL8/KGbKpERG0EiB2Ro0ZIisQuAICYpZSIqCgKRDQwaaJQZGrM3CRFaOw1kIgcc2eLhEj9wdC5XA3M46NZ1o9C8B7y0wMMsElmKCLUDJQcYwQAYgcAQIBEIrIpyxxnHY3H/X6PnIsxppTUjIlEJaWU73tq3fwBMedNzA7SqiaZmFQlaqKlaiYiSSISBufz8CAimvJI7dUgiSiA96HfHyhiduYRBVS4M3I/+eDtN87Pvvve45/96vOPP/3888v51XxTK7S3urUq92+9p/3LRl3X8/l8vd4MhoPRaLRYLcuy1M4RaytBBshdmUDVkiRQJKIuWNI9m/N2jRFUdxvC7iewG00kAsgm0WZf8tRUg0pgWcnldH7gLPQZCFzgQfCEaKrDuhYDbWLeZmA5pIlN3mkQNbWUBERltVTRyIyeuSh88K4IruiFIvgQgpFHdVauc7qGlS+d8Kurtccee+yxxx8dewJ6jz322OPbB0a8hOMTTwRarZfValZvlrFOeY6aYsxLhgEMwbJJsWMCU2IPJr1+LxSFCx4wC5IKdAFcUEfZilIlWlSLSWO9WZfT6XIt/PTxs6ur6aasoZ1Q3JK6MNPBwWQw6KtqWdUxaSj6VVXlmXAHInbO207CwMziqUpKaGZZ1NXqPW/kZOvY5zytZXZqjReBYwcAkkSSpJR+N2Ee3v6jI9DAFE1RMxcB2TyjJVfBlAjNuKF3W6sMbGvzMgHdyU5h1wmjIWwJMhvb5iJs+efMHzbKo8yAtEvOW+a4JaM7RVEm9Vpetd2kmb21fF4jrstLaDM3rTuFtax7R0/fYBCb+mdKeuub0LEy2aUEttRzLqfhorFxHM5+1NoR0NnKJEWRPhM5kuV8FtgPJ4jshgcnp/fScnYZy41qObu6rMpqMByH3uD8/qOLF3R1dX3x4tlqszk8PLxzfHp4dKeuqvn0enp1oej9YHJ8NFHVVMCbZ+OnV4tPL6ZAreE4ADOrmookkUwkiSQRaU+nmZAzkajma5Vp4o6P3iFwX6ZOspeHmJqBcqaJTfNOIgKATBRTVFUEJCYAFEn5riUiFanqGjGz3m5HlW5m5usaAZNE5xwRdzrk5p5CbG2gd7JrQtcu2RkgtwtgEx/QnfPIT4C2dTNhlUMLaKaGBkgIbW5Ma0nt1gUBGneNpvO1USho3J1b6w3bBoR2KOpWVt/5zWRvBBXNzaUq4ohOjsb/8d/8+Y8/fOvenYMBGxM5qVaX0+nl5XpT3j2/Nzw6MbXNfLZezJ33k8PjYX9osVrPLlO1nk0vylifnN+fvPnh+PRsNZtePP7k8snTXn949vANP5zg/EV3f/xJwl4P9hlgd40LAoKiAYExgCfsD4rJsH80GvzZD9754Qdvf/jum+fH41Gg1fRiPbu4WF73HTGoSt0riqIovO+J90mSZ5+Ndwof2sRrQETsPTFnYxkzUzP2TNS5UJNjB4gKllJCwuBDFvtj49oPkhIRO+8pxZRERABz8kCfVcwpCZgxcfCBHZtKDjbGlFQMAZVZVauyRELvvQ8MgKISY0VEREXOOJBSrTmHqDRQQHYueK+SUqo3ZZlEzIyZU4p1VedwDxExto9sAjPLKRwAQLPRjYFzzMRN2SpqxkzRNRRhrJOpoKEPmYBWZEw59TGYmNR1ZUDE3vvB+dHwwdnp8cHw3snweIS/+qz49Nns+Wy1qqROpgDaWn7tOejfBSmlzWZTlmWv3xsOh+uylCak2sWbUW3X9MRULaWUv+V0CTa37HMXw94S0NsvMu0QYK2hv3nHhNAGccnglVpjBABRK2u5mi5OenRQjDEKgTrCvKjIhSIws/ecvc5ANYmp5BU9pqKSlfqKoKox1ZtkGhFj5ULwtfdV5UPwzntDR6HyldRllFSjDeve8KOPPvroo4/+MI2wxx577LHH18CegN5jjz32+PaRyAdfOutXq9li/iSuppai874oCnJ+U2pVStJU9AfOeUD0RT+LNJ2ZI+oNer7f4yIAGKiiCYjoZpXm1xKT1cmSpCrGsk6itZgIzFbp2dOns9mmrmSrfOyI1caCgw8PD/r9XlVVZVlXVc2G0OZM75Bp0zyTyfIrEcna0rquW0mmddRqS7CCGYhEEUEE51xd14hgYJIEAMwsxrhaLauqkq0C+utPVjsaAZtFybidi2V7DWglzw1Fmpk4x9ysPdZW5WpoitaQmYCI2k7RGn10Zt4QoLMc6IR8DcObZaddDreGee7o4BvsXnPUhiVuymgdMDKv1zC/OwR0Z5axlbu2/GOnckLoTrmTxSK8dOi2yaxJLdfKwBvnaqauUHwZQAaturVhc7NfCRIgWYz12PnQ7zuI8/VqqQa9wTgMJ6fnb/jQm18+j+VmtZiWm5WqHBfno/FBWa3XZbVcrTb/P3tv1ixJcp2JncXdI3K9e61dXQ00gAZIgBSXoTgaycQnmelfzE/h39DbmP6CnvSoB5mMNjSNoBkKHBBLr9VdVbfq3ptbRLj7OUcPHhGZtxvEACTAJgf5WXfVrcybsfkJj/TvfOc72xVoXs6W1WR2cnaZc961jd69WRLWk/nl5Wlj228/Wr54dfv67eqmid6H3nrDjIicYxHNOccY+wuCVDjQqgqqFmNkx8U6U0TUFBFEVESrEAAgSzYDIgrBFxVzTMnMGKn0d+pi9N5770vqBcycYzOLMceUwcx7F7tcTKWdQ1WTXJItUshZ5t4bWkWZ2XuXYt8JqpNkFnti2HSgDwwGgT8TIxZqG6lkNQCgWDsP1s8IB8mM4d5EtDEeykCXuNDeP2TUKQ/yeaT9XVnyFL20eXBd6SPHYNylDVmRQ+Z7TE+MwVNUmr0KWglsvpz9wQfv/fHvf+O9p1eni4pyp7lbvfzk9vY2JpmfnC8fPASz7c3NZnWTcjq7uFgsl2jabtbddt0122w4O3tw/uTdxePH2/X69Yc/ffXiExF49t63zh4+bmPumt16ve4lqf8oEfQR/zAc8M6AMBQugBmhsUGFsAz8nedXv//d9/7w+x98890nlyczlDbefvFyt0KNDHo6n8wmtXcsplVVBRcQycRMLTiPCKbGjkuuqNwUxAxICiCiAEaIRphUU0rOOWZqUmJm5zyiqWgjXdM2OWfHrqoqYl7d3RHRdDZLMeWcRKXY8k4nU8m562JfhAHGiJZhu9mUey7GqKoIRISFTAwh+OCb7QoRVWS9WTvn5oslI5pBFi3tEAgxxdjGThXY+bquU+5STmKKfaYUc84pJ8eekBBKY4a+4QEAxKZJKarmnLNzbjadOSKz1DQ7My3pUjBHxKqqWSTmEEIIvmhgHSAi55je3t05x0ggmgDJkEW3QHfsqhnidx4tTsM3v/vuow8/v/73/+/ffvRy82ZtgpCGR9kR/0iYWYxRRKqqQoSYesvv/iuNoWrE8d9gZiClVcRIQPddAe5hmOHh8JZkoqGSBY3MzJzjkl81ZRNRQfvytNl/3WAwFL1brVdz1yzqTbOC1HlC9uw8B/azyXQ+nU/qqq5DXU8cExMQmkkSSSJZJZuKc4RkAEW6byJSHjCqtlu3XVw1KSmwm8wat8hdslnozr4Hu09/m4NwxBFHHHHEr4ojAX3EEUcc8TXjh//7/6pkqN5VlaS23W652DoH5z0757z3MjMxdFVNyKrqfUXs1MxEwAwdi0Buo6SUUyexsxwtJ80JVUEMRE1MRXdt22aLFD77/PqnP/9ws2vNzBHYLxKuFAKa2b15c7Ner7e7hrMh2pfKMomY2RfhMwDknIsCGmCvi2EmER01mIdv5ZwLiUbUu18WYVfhsptdm1O2fzD7PAJx4IbLv5CQBr4YCw9cBJ+DBUEhWHvhc6/zHHnqvW+BjZvfa5/RgADM7smKAAD6HlZmNDDDg2HHQBX3BPW94z7k6gCwWD/3NtbDmeHB7w8OGrZXN1tJTRTCcfDwgP2mRwfefh+jpBUMafhjGILhv1ESDWXTPQ1N/V5Hz4XSvL7/dQQwNDBwLsxmy9ly4jpKzd1mfaOm4KeL03Nmz+hWb19uV2+wsxB8N1+4KvhQn51f1XXdNpu2bd9cvz49PZufnKN3X7z6bLu9Vcsn5w+m84uTuXz74fLuG1dttr/55DYpEDONiRPrzxERU0qq2uvPiZxzqhqqwMRlWV56lBFRziKSHbvyepaMgD0BbeZiBIOi3jKDelKPunIiLG6wIgIQnXdDssHMDKl3sMkps+O6rg2ACIMPWSRnV0rjx9IBd2APAmAlnXKYBoDi9z0wCINZB5QBMgMthph9MIyf1tI+sI/1IT0BQ3JEQXXIXpQem4fiONwH6yBwRkQDMxoiCcbfxPFmLLz4cBDlyPu9FkIcREDAbOL5+aOzv/hvf/+9x2en88qzdZtts7558+rFbtecXD5+9OQpsO/evt7eXXfdLoT6/OoSsjbru3a7k5yy2vLq6eLB4+liGVc3r3/+8+sXn0jszh48vnr6Djjf3tzcvn558/Z6SDj9DtJjv20tKn71J7sfG/cvuyEYKbLZog7vPr58/ujy3YeX7z49f/Lw9NHlyUkQnzcW2wDRB2T0jtAzMe/tlxUA1UxBs227Bkpy0TtAyKXXbdkx9m0DAdDQsoiaEXGX2lJ85J3zLpenG4CVeQMUSimDqoAVjyxRkTKhqmrTNIUjy5IRwDHe3t6YiubyUOtdzsvNW2pNcs5mkiLknFOKXdc551UFEVU0pYQAhBS8zyIxZgNkFQBpdrsudgJaui+oWlExC6AY5JQIyTkOoaJSKoHomDOYc1ga8CIREy3cIouoSumeq34TphUAACAASURBVGZd14FCPZmEUDFR07QA6EPlgsuSVTOCAZrjQMxIzsAZOCQEszDhyYOTi5PF5el8VvtPrjcv3jQffvbF69vtqhUdHkg2ZsR+1UD6Xbs9x0fyAazPgMfYpZSm01kpuxGTfsInxn1qcsjuFZnCYP5VEjCjFdXB/rBvZzG+gjh0me5dpNTAOabyWFc2ZlM1ta/kFpCAEETNdl3MQNPFCVUOpSXNVppOAKQUN+tVbLjxLgTnHFfB1ZVnAiIIwRG60t3TETnHCFRurpSlWIDkLCnFaUqCiN57rjukNQZ481fIF7/5MTniiCOOOOLXx5GAPuKII474mpGBnKgF590EcwOAvqqrQD54JnaOfajQeWAH5FU1d5HIETskkpRyjJpSSjmlLqeYuja2jWoGUzIlREZCIEeO61pTTjm1op++fP13H32666IhEAKNFOGA8gX+9PTMOX/95s16s921LQtwEVONbe0BnPMhUEq5KC5HJrqY7cLAguUsAFacnYu6ufB9RTGtKo4dO8eMIiJZSoOd2EWR/NWL9qsA4YB0xp4fLcfDRQk2aH/pYDGGgygYkMAUELjog0oxNhbFd9kkDE7M0Jsg9HrQUXJqeMC5jLYb4xUehc8weA+oqJqq6UiEDyfSs4K93pp6NXWhggf6uhA4ZkOn+z2JCGVhqKbSK1X3hzFcrcMjHC/b0G3SBg+FQbnd+36Agaj0QtdROTtsxxDACAjMgEajDgJSqEO1mJ8sThbprmt3d91uG7NimBNxXVdnl1dMcHdz7R3tdpv8xaenKbKfTKpZcEwgN2/e7ja7GLvLhw9nJ6enkn72dz/a7LaK7MLsweUJiBg9pXpxvf3bN+vsqqqe1MwsWWKMhaNCoq5rc85MXICIasXKtI+VMc6LC7SZERWz11Tq3Msl18mknHKWXNylc84ltp1z3nnE/q3gfcm79EmP4YJ1XYeAVVWVlmjFBmSoFSi+tI4AvXMiWURxHBnobU5wMIApXiulv1nfe3CfPxj0xkM24hADF7RnLMo+VKWEpQ2JhoOQvme8UhTUYx5nv9+DpM2gze8V0XBvWyXD05+yY4kpIujDy+Wffv8bf/Fnv/fswemEoN2sV7c30m532+3J6emDx4+pCu3rl69evpAcF/P5+eWlma5WN3m3A1U1OLt6OHv8rpsu4nZ7/fLFi48/ZrJ3333+7Fvfhvm0ff3mxc9/+slHP++69n4G6HcQv1Uaup/Q+qkK4CuM83gEhmCMEBiWVf3Og7M//6Pv/MF3v/md954t554tdbu1NXftLjuwOnBVVwhAAGCQJYsII8WSXgKybDlJbFszJUIXHGDxZ0cAENHesNl5JDKEmBIgTiaTruti7IL3KiI5S/GlBSAAIgIzzdkEGREJTTKaEYKVdwHbtsXB6wARmN16tc4p1sGXOdM5p2rlSBCR2alZSmImbdd2XQuA2ts2mYjklIjQscuhMkQxQyQ0zZK7FLsYBdR7X6YBIiZERBaRrEoIqIw9zw6hrs0si5RiDnaOvfMhVHWVUuq6rlRZtW0Ua5Foulh4H1QNUiakqq59FQyEPecUwdQ5ZnbMjsgDkKimrhXCWV0vF3x2ury8OL/etJ+9Wf3Vf6Aff/jFi+umiSlmzb35y742aTAJ+vtC6Bexsf/146tnXdwysG3brovFhdw5Z6raJ6uL/cpB3RKhAWgxRiNiJCRk53LKYge3fl/wNH7zsXETAGCDVxhasaiCwUiMgAmMAL7EZZcnAWbTbZQEXM8Xc55WmEA6kZRzVhHpUu46abVFQwTnuKr8bFr74EJwVR2C90RciHXPlXMOiVQtZRFRJEZAA8siCgYEd+ZtknZ3mRtn9Oa3P0BHHHHEEUf8l3EkoI844ogjvn504OsQ6umCK6sr9gGdAzQBSVhY3RglN8wsSdqmkZwBIASvojmm2HVFAhOquvj5eRfIOSxlxYAcaj9bLJbLucjN3frnn7y63snnN9udWIKylgAEw4EPMAMf3GIxvbi89M7tmlciCqUfDOLgqWAAJiIpqYjFGAvnBQAAmFIsDq5MhEiq1ityQa1XOxqYluaKjBBCAEQwzVGhCG1Mo8hmsxl0aoe0iH1l8Ym/gDfBsoIiA7C+hSCTYxyEx1wawDOXpdXgj4nMTIhWVLwIXJwzy3VBREArYtDSqsdskD/jyOLuFcl7qfHAugyk8qEqqV/XgamYjWdnh6cCRch8wO0dOhvcx+BmQPtj2lOMhwzkaPkLB1s+WPfj/au+943GYS1cWO1x63Coi8bDz+O+IRIi5AQIMUdyPF0sLbeSZLfZ5vxRu7w5Pb+YzZcnZ2fvvv/BzfXLZrfJ+VYlz06uLq4eEU+zyHyxzl27vbsGk/NHT68ePN7uVm/fXq/WN4D+4YMny5k/6dLpRJ8/WK7bt4BIyESsZIXizJKlEyQMITBTzhJjrOvakcuWRUQBSt09EXZd6z2HMGnbVlUBtK4rREwpFVuP+Xymql0bC61c13Wp3y8rc0DMOVcuzGZTM1BRJKyqyjufRUwVTAmQCIt0sYxQsYBxxDnnLkbvnSNGxMKDY7kTRXpf78HHExFK7z4Y1NHj3TAqjQdnjEF4XF7rBf9YblXs2bzx3UH4puNGx8zIl7IsB8M+hNIgfB5+gEEsPUTSEJNWPHBUNEs2M8o0qfh777/zb/70986mOmGBbIzsw+TDjz5ZnDw4eff59Pws3l6/fvEZEJ+eP5jPZrFtu3YLElW6Lnbop5OrJy6E5u7t25df3Fy/IaLH7z1/+OwZTKZwe/3Rj/9mt11dPrh6+k7LP3oJWeGr5/Bl/H1E7W9bR/zPDV+djb+KMuKl5mTMCpaJedTIlwSIMQIBEAAbLCv36Hz6Jz/44I9//9vf/eaTs3lVu4zSgYlzCoqqoClr1mTUP4pUDVBUU845JzAIzuesKlpXFQJ0MTVtkUgGXwViKk4vliTn7LwPdTWbTgqd5x1JHYjQETt27BgMNOdRuVxSJUhUbGrZOQTrckI2BLIsokUmTcyO2VeTiWNmopJnct5j8dboNdGoOYuCKpKrJ64udgqGkFMyQF/XTIhEAsiOg3dFqc3e1cRBlB37EIIPwQdDFFPJYmYLAAAk4ioELo7zpQiJhkcjO+SiHidW8VmQ0NQmWarZUtX8dBJCRUR+OgMA6q1LLExnqqnovsu8wOiKgbv33pmWNOmE8Oq0Pj+dvvvo7On5/Mcffv6f/u6TH/3kxWevV42AAAqQDXU1vdewyL0ww/sZCgCA0S3nN3jT/Spbs18t7P+xezzYh/2iMy0/63azns9n3lMVvHeua9ssAmaxMwQAooOvDcVtCxExZ1RRQiraflXF0qPBIMdIxC5UKtrbnRMRYjQrSXCVvkFCzghYciNZJO/d/Ie0Z+GwFRRAO4O7zt5s4+vNZno2rSeVMwSo++dBVsiiWVSLt7mJahvTpm3VFNCIkImC93UIVQh1VYcQ2Lk6VCFMsE+MYyi9ckGAJ7nGT1bXaJ3l37Vp+YgjjjjinymOBPQRRxxxxNcMQySUUFUuOG+1QWI2gCw5SoyaIqimLqYuFh1Wu2s0C5h1hRk1kJwtJRMB79l5DBWHwL5i543ZnOPpoppMQ12DSgvev9012W43bVJQIDMtzE9hoAvXOpnUy+UihCBqMeUQJvO541ATFNYrFRpS+1pOZiZVY+bBoaJvleTY4YHnRmGoDSxnYaLgXNdFM/PeA4CItF3rnQ8hmFkRkH7Fx+JXxJ7y2BOiA++hYGiAaGCKikCIAoNvCACAYlGBFrJsEDKPfRp7LwLCPSFbrCcORESDSJQOKOeDY7OBjBt8dMEQgHiUk375ZOxg/8Na9CtXpucgAWGkn4uUDBEHYbaNTQUPiOL9QdrYFerLxzEQzzjobIvWuphBwoGBNB5sdGTAD4ltAhKJ69XtbjM9rWm5PHWE3vFuu9qtsmdgsmoyPb96CIj2+otmu2p2G6JqHarpdDqpp48fPX7z6ouuaXPs2u1uMpk8fPCYme9uV81mdcd+eXJ2dTp757J7MMdlhZusKcUsNFC3fYM7h664JKuqqKScaPA0H/hcVAVVJUJVNStSyFzUZKpS1Is5O1MoSRcYjGgAkJAMTEUlZ3BMxDnn4ulRLmGxOrbSCLE/ksKHWW/NISJSWpZBYfuLkm1QnYNpiSKyoZtYafxXSIDB0sXGABn1+bhnpw/GHMCgEBYEJaJBDUrvwmLHYrDXKh6YhB5w0mOMlqHHg/6mB5x4OXobj6rYz5ToVFXJOedMqL//7ff+/I8++N43H12cTlGiZOnauNslXy0evPON6XzZbHbrVy9j25w/fqeqJzlnEAO11e1ts9uEavLg8RO/PG3Xt28//+z61StVePrOs4unz3gy3d3d7a6vg8nF1cWK59XkGr56+/0a+JdNc/yiOeU3uO3yFx68dG9yL7X8DBAIpoGePXzw3pOr95+df+8b73zj6dXZFJ3udNeJZFNFsNKdzFQ1UUTIKauKqZUHU5acs5Q9MrH31WQyQUSR3kudnfPBIxG7hIhMXKpj2Lni2IOESMhMpqpqUaNTR0MKtpeZ9vcTIjGCEZEBMAAhA6ALoUwIvqqcY0SaMReWvBxGFQIxA2DO/YQjkovDDjExEQCWWqKUEiLWVd3rWhFLPQ57RiQwq0QQwTsPUAqYgkE/Y/QTWUnCMTt2xNQXypQZGgmRDHt5LDGTKxbzxs6AWFWZCZiByNc1wP4uZiayfvIpKSoCNhASQe5TsqhKCsGTDzU5XzPUDmeVW9T1Tz5+/fHr29tt3EY1AyNEIoU+03UfIwO7z2v+RkP018I/A/318BROMXZtm2Jk5jpUW9gUIr84tzj6UvK+JLzRyuMCDQVhaGhMgEBYsvIDh4yI0DewFbWxTQCAmUnOVu5cQgYSs96gCQ7T6H19nRg0Am83zYtXb+aYnPgas3PsHDtidq5U+SCCARbJf4xRNGcV0ayqphqzicQu5l0bHTMRVSFUIRCjY3aekZlK3+hJFcJUVbIaVPNjH8IjjjjiiH8OOBLQRxxxxBFfN8gIyLFjz5QhSbaUJDVds05dl3M0yV3bprab1BMw6NqWENBAszjvg/dlwewU0Hv2oQo1heB8FeraVTVPJnByYga2awGUHNfTmQBsmq5UKioAQuk0B6NGdzqdnpycqlrXpSw6nc/DzIVqIhIlR1UpBhow8Jm9JyYUdw7wngGg+AYgoqmWX/DeExEg5Czeucr73a4RkbLgyZIBoK6r2WxWehgWj4Jf/5oesM8HMFOVgaRFVCVEROp9QsZzH8yCjQdfjvLG4H+BCEBEpdXb4OLcF6oe6CYHKfSgbu5X1KMQuOyOCPWAkem3digzHt4yMxzIxJHrPdgX9BLtcSf3SL9Bg9yLWeFQ6Wz3/hopxfEA+hMnGuyBh731bh69PMv2Hy9EZE9e9hvfnzgSgea4W93eXfPsYj6b1OHsIjjOaZdiu1m9UUuzk9PTswfTxVJEiNxuu2l3GwSDfLI4Obk4vzCR25vbGPP29sYkL8+Xp4sz7fTu5u7u7bV3vp6dPFpO3j2rPp679jZvdkkNnHNVVacUBxYYzTTFVDjfpmlGZ5gi/UopIQIRpKQxJlUpZtAimYjNNGcpzcSKN0uRgHVdx8REZFrI56yiThwhxRjVlJm7GCHGnEVyVpUqVOBYYu9+bgBVVbHj3W5rao6diBTC2nvPhCllACtOAoTEQ9u+8mtDxsRUdNAXD0r1sbfb4RAPmYXhp4PIh0It7fmgMsLjiI5S+mGD+yTJECX7oYchdvsQtEGTbVo8cHVIiGkWUH364PS/++Pv/avvv//obBrINrd3mi1lQApP3n1/MV92m83m5k3abRfLxWwySSmmrq1DyClv2wjoZmcXiwcP2rZ9+/Ll7fVrlXx2+ejBs2fVbLpdr28++yyuVqdnpylM4U1smuY+Kfqr4KsT1AEB8y8H+HUcN+4jwxjNEaDiPODDE/8//PEHf/qH3/vuN59SbvLu7vbVFyCJccihqKkIIharmYEK7o+d+rQoIhH7sJjPZ7NZKSAAxGJSkVVgSI4654L3hCiqXYo2yLORGQFz7mLXxZgIC5ftilVSf8MgAhI78o4LtV1XXGZZV2HJEk0nU0RMOXvvESCllFIy06qqB7Kv3M3Yh38pzyF23knObdeJqCOe1JPSe9YF36XYpTRfzAGgaRoAICLHLqeUUyrXggBc6JO7zK70kCiGG8456C04zAwUoLDqpsLsHHPxVgIA772ZmWnOyQwK64dQKi0EBqYYAYjQAEEBEYkZyUp+2rrONDPixIMPuGF9dFLPJs+uLs4eP3z5V//Pj3/2+U283ZoZIAOBZTG1L99Z9+KyvEW/USXyvzQMRiWqklLcbraMOJnUxMxmSARgxS78/ocQgLXvBd1fOudcmeyJCJHAe1UTMWBChOIODgAZEfqbi6R868sGaOwDI4BqtJhVvzRQNmTGDSAD3G6bjz97OdVGt2HmtK5CFSrvXHA+eD+pah+CC3743lWmCM2SU06569qmSV0UkbhrJGfVPp/kPYfgq8q7UPngfXDOfAohx06y8vMfrNf/+Z9gTI444ogjjvjlOBLQRxxxxBFfJ/76r/8X3GRR1tisXm45rrW9Bc0mMcWuiKQY2SGbrwzIANBXIoZEYVIRMTofJhNy3gCByHnv65q8R+eIgEysWcfN7Xq1url+M18suwx3r263N3dp25qMBNBov9ETtyfL5dXlVdulN29vXr16rTQxCjEJgg7uFFZkWWbAzIO4ds+EFjJMVZEI+4UNxtJDich5b2q7XTOIScnMCGk6nRY/hK5rm92ua1sR+bWEToMnAMLgM2CI0PsPQM+jWZGTau9Xi4MJRSETTAonL8yDSe8hGWyFd6aefEbaG3AcclfWy5x7DfDe/mIQFh14Jg8yod5KsYhP9zvFUSPaX+Wx0PVwb78Yo69Czy+Nmxk+ZIMBQyGJx96FI309sMu9YPvg0A75qj0BbfdVzzh4TtvoQ1IzSE7S7tbXuqUY6KKezaaLk8lqBpC7dhtTmyURIvvJ8vSirhZfvPis3d7gNgXWOnBdnV9ePRVx19evt6u79d1Nzo8n0+mkmjVu227bu7c3s2xz9t9/9+LDl7efXq93G8lmSES02acJRqJWVc16yTti6ZlZ5IdgFjwX7XMxfVZVQGQi772q5tzroIl4lHoX7X/vhmHgnDOzm9sbhLHdF5pZTNnMCKFtuyIsLwwys2u61gAkpyLhLHXNhT8qPhv95S5VCEWnaUWYOZC+poXSHcJvzwXssyoHGYdBD3n/bTAofSSxj+jxA0Moj4rqvUp+fzsOovqiazuM/738eoy1wmmpqimazSv/Zz/49r/5b77z3XcfTFxavX179+aWKExmZ+dnF/OL85sXH928/lxSd7KcP3j4MLed7HaqIoTbXRNmJ6enp+dXVxHs5ccf3rz4DM2uHj5+8t77OJ126/XdZ5++/fzz09l86ievN831Zy/fXN8U6fr9bNJ4Lnbw8983KX1JRvwvWxP9G0UZdBmu3niFS0dVcwYz4icP5x88f/T9bz17enU+x+7uxUdoUXOXYgMqhFAsjwhR1YjQE4uqmTI771zxvWFm5z0zlS6+PgTHrEVZTIzeA4BlgyL7JVOiDGSiIpqNABGIigiawMiFqp4Psz0x85DLKWeFBuacCyGoCiCy86UUgZmh+AGAqRqpUUlbqnpRAKuqqpgemEG5ewEUCZ13ZdpXVa6qxXShBgTASGpiZuTYERt7NQQA5yso2VMk5xGJdZgWilu/eSAiVcttW+SvWDogSuorJkSdYyRMIiiqmiR2Ztb35u2ltrlMggoIxWxXREUOWWAzyElizl2KzrsiCd+uN13TEHFVV+zc9dvb9a5rkwmEByfhT7///OmTi09f3/7s0y/eruMu5cGDmBH0/lQxRtJ4A44s6u8cEz3IkLWkp1W1nkzZ+V3Tln4DvUPU/Uy2AYxpeDVPSOxYpbd1GpPfOHZtOCheCiGUhwwxe4AqBDUBROcdmGpOiAimUdJXj7Y8rhyAijZtbjvdNpK0ZWwdEbuigPbeuVD5SV1Xla+Dq7zzwXnvqsrVNcPU23xiWUrupFQL5ZyTZFMVy1klNjvbAQDSFmKdcicK8PLF/3ZWf/O3ORpHHHHEEUf8SjgS0EccccQRXyua2uatu61JY7faYLrDtENLVrjhUlDsnfOBXb/oYiQDYueqaoLIRFxPZ8SuaMJKMyUgEs05Re1abXepaXaru93NrZPcCN1ev96tNhJlWMX1vg2HEtjlYn5+ftbFdHu3urtb+QmRR41CZIRWbJOhF15hMdAo7gFlYcOOTFVEiAgA1Mw7BwAp52IkEUIAA+mdB3tb27ICTwnMtG3bpmmKiec/DAci4cJ0UGkaP5yp9SsuogMOrDClNgiLFIAG9+pei2Om5aXesQSBeo9FPGBhC/FtA5+31wCZmengXFnqXQ8+V3jJ/e7uGTP3HHRPQO9Z8ftC6f26dOCOEQGBkMYzgDIkMDLbMGy757UHOr1cxr5Dpe09qHFcpB7u3Q7/HzEcyaAWB0PELKA2qWtC3KzunGP2bjafPH7ybLterFY32912t10n0ZPTy5Pl5XyxvLxIL3Z3Kmm3WUuSZtctzh7O5qdEvF3fvnl7/fbV65OTs/l88fDB49evXqfY5Wa3PD39vedXL252H1/v3m7vYoegli0776D4rg6XrAyBY1a1nBOWuNXe/sIciWhKqWjWAaCs2IsIuhA4oCZiA0UP2XJJ0hAhswOALNI0jXPOMROVQFBRRQQjEk0AgGhjxqUsr9EAEQV7VlRFcRBeHlzj3nWz74pZhq1X3A9hc3BfjIxzL3fufxqSDIgDpzxkpsCw555h0N31MVZswMsvj8ExKqrH8BiSFuPB3JMZ41D8DeUMVUXyvA7ffv7kf/4f/+z733p6NnNx27z84jqwXyxPlidnoaq6m+ub69cEePbwwdnFicWua9feMYO/uVs5H66ePZ9O6vbu5vOffPjzn/5kMZm+8943Hj1/j5Da1d0nP/vJzauXs7p+9OixKXS7drvZ3q02v1QA/SVy+b+II/tcsJ+KB738GBhQoosBzhbTZ5fL7zy/+O7zxx88f+JBOG3bNiFpSSeWhBAVoW/wKkpErqrZDACCDz6E4D0SOcc+hNKTLQRfTF0GTpZLvpORgAiG3CchSU4AxIzEhI6RuQ92Jw7ZOS60KBGLFZt1MCAANCy9STmrIKBzTntOnIo9rmoGKk3dyJCYPbICALADRDNDJFLVLH3bYOTeJkiMGIjYM4OZ5IxIRCWBSYRULJaZWE3BTFQQgJAUFMqdNQR0TimnnLrOHJOppFjchKzsSSR4T0yxa8v00rUdmDnX8/sAoCIqOjzEtG84bAoHM5EaZNUkkkRseFS02yZ1kR1nyeycSCLUwDCp3HIxu7o6fb5LL282Dy+XP/vszSdf3N1s2jYXlhv3VTRfDqkxiuxLXe9+V3BwXXKW7XZbT6b1ZFJVFUYEMBuSLofAPimPBlDc/glRh/x3GVkovamBx0x0n7zpLziq2pA9pz7Xr/d31T9Z771Q3s5Jt7vUJcjKzjwCZIGshlnQAWJyXdw2bRVcHbiu/KQKdeXrOoTgPJOrPIWAMKQmzFLOKaecU8yxSzFnkaQ5a25jp61HYrAn8KTrbn/jI3DEEUccccSviyMBfcQRRxzxtcIc3Jy5kIIjiwJmnllNGTn40HVdzpmdd84Te7OydK2q6dSHCpnBEJDQB1O1LiaxnFMTdzl1KbWpa1LbSNc6U0Y8W85DFbar9ubNTdu0A0H6Fd0QAhHMppOT5fLm7m6z27Vd5JCRVExTzGa5cLJmpfegMbsiyYwxigiAlfbqRfWcJXddV4WqiEChl/CqYxec67rOzIqbh6qmVMxzQVXbrrvP6v5qV3RU4iIVZRBA4T2074iDgz+xGSKi41HB3Gt/Cw/H0NMNfS/4csrQ68yKJcboRgED2wsDmz1QbiPvNkiDbWykRP3qb5QCIhET7s95NJnuOdxyHAbAVoTX94YNAcoSEbEYJPQMyWivsP/9gWA84Ir7Tfd9Fvf08yCf1Z6V75nFPQd9QG3CIKdWU+111eXUAYs0uvAh5Hg6m52cXYZpjGl1e/sma5fzWQh1PT/PELLdrte327fXJsJGy8XFyekJ6vPt5u12s75b3TVJuFosTs6qSc0hNEna7brZrZ3j5fn5e++fbG9v7m7evn65np+e/uBbT940oPTp335206kzs7quVXWz2ZRKd0Ao/FFVVSnnZtfUdY2EfXgTTad1zrnrur5lJaL0kjEyM+/NOZezxJhLeTIxqaiIAEBVVXVdGQCnZKbeO2bHxDHGnHOho5FIRAGAGVNKxcfWkWMqBIypyphuKE6uznGxAilerYXIHry/EQCgVyYOWYH72YKBIT7MKAD2LcnwYDBHXbyNuvg969NTUQYjU71Pi+C+FmGI5OF27vMiJUxLMJUsjqp0MZqZR3j30YP/6b//V+8/OZsHNJEsVE3Ozi8up5MJgmzXL+/ubn1VLc/P54ta0+b69Yva+Rht10lE9+iddybTanvz9vOf//TjD3+6WCzeee/9y0dPiJw124/+8/93c3tX1dPzh4/c4sRijOnVdrPKsbVfzEB/iUq2X/Ti4VtHfAn2pZ8RirZWAYzAHMA3n1396z/81vtPr04C5t2dSXKowROjY8fkvJqpKSJUVTWfz7IoEdZV5Zxjdj547xyzMzMiKj4bzFw6gqaUqtoXX/WUk6pyKLRzmYWJ+p6ivWM0OWeEWUSzkFMmcuy0ON4yacpggIxMDomBUES6mNQUELJKuTfAJHVtjJ1jLtpnMyRkF4KIlJ4HCEiIzIxWvOYJELumzZJUpRi+dw1O6gmC7Zq2CsF7V5I0vXsVESJqTpKzihSLDInRzBKiYzazmHPbNDklx6zOiH9LsgAAIABJREFUZabYdSJiAFaaMIo4dojQNg078s61bWcA3ru2aUWk5EbNIHVdbxNkRoTOub39T8nZek/sDHGz24hoVVWOeDqf1SG44J33p+engGxGimTkiOuM3Ar+yR/94Ic/+un/+e//43/68eevb7eGqjbWXwDcL7kZ5hYCGEsWfrdgWpo0Ihh0bfv69evpfDH3Xk3btikPr7/no1g810SVEJ3jLFKUBCqSZWhgQI6pv0NKVUrRUxenmvLtSDSLCgwPezTVLGB00B/y3hcEBWhTXm0sCfpqejo5qbxjhJSSghmBWZacuy7uthsEDZ4qz3XlZrPZfDqZTerK+f6RyaVjJnlmDk61qk3FxBQka4qpNd9gtVTWmMU7luk/waAcccQRRxzxy3EkoI844ogjvlakAA79ZEqOsgtMM3ZTj+aIgveViKoSMzIVSSaoWspkWZNap6amWbqUcoqaExGaaspxpIbIBB1NfA1ASYCqqbKtmtgmGdUq1Atm+8UKE01rv1jMp7Pp51+83O2aLNZ2kQTVEEAOil6LZAZUpTBxOJppUG+fbGCE5H04aGsDWFo9MTvnyuK39Fgn4iJVyzl3McYY/7GXt6jFRuMIJmIuKk8aDDDIuZ6AHrr24cD7qgoAMLv7ek2jPXfWf27kf0flT+GeR2p7rwbuf0CEvrP8nhdGpNK2aVB3DVJXHITF/S4MgJDutfMavRP6D41a2PFjh4pqw2K/C3u98uFVA4DR43cgkXsu8nBzPaM4fmTPOKuq9FXqCsMFGcTcZjXZZDqfn5yen2NaQ7d9u757a5pPzh9OZsvZsjL0CsgbyV23evvGEiyX56GeIF2oYby7bdp2dXdrRmEycWFydnHZVrxdr7abVZhMTk7OvHOS03a7QqZ3vvH4j779+HrV3u3iF2stNhxItFwuC/NqasTEzITESDzFUFWI6JkHpbmWWv7xQhXn2ZQSABS2K2cpNhpMTEwppkIPERMRqSohhRCGMeydVUWH9oP9ZdYQgilkyWBGgOycgQ1898D694t/YZGRQDYVACs1B1DSAPuQHKJuEDoPyZGDomtCQu6pYBg01QCDWc09ArpsWXUfzwdx03/6gJ/Fg3RML6nutzaUEZRURk4JAHKMJ/PZ97759M//6IPLRYDU7VrJ2c4uHi7Oz3Nsduvb2Nw4B9Pzi+nixHK7Xt0RY8pxt2sF/emjh5Ozk3h7e/3i4zevXtR1eOe99y4ePGT2m9ubN59+dPvm1fLk/PLRk/nyVFTfvLm+uX2DoBfnp/TRHchvSlB5cLv8C8LeEuU3sbH+T+v7ovY2LAqgCOYAFlO+Op2/9/TRd54/fPfq5LTmisyUmdETVI699+ycIpJjcpxFnGPwVV0753xVBee9YyYmMNCiJmYm78sk38Xi2w6hcoYUs6QkBka9wzOJKmjunYKIiChK1pwEFMzQwCNpyl3TqAoA9vUL422F4Ly34tGjGRHIsZlplq7dFSstrmp0johFTJHUcupiSgkJS00LFRcFEedd6eWrOeech63K1rmS8fXeO8eF7zW1qq4MLMVIhMWM3rEjohRjsQEpKWFE7p8+asVdGsByzinGkmVF4l3OfedPJnYsYoUlZ+bgfRUqVRXNAOhc8L4CGh9xfcCoqSEgO2JCwul0UpJws9lsOp2WlAAAhKoidoCUxBSQOGTDZHBhNK35wcXy/fc+/eGPPvrh3/wsgwrCQSfisX6ipHtHD+jfOfb5AAgAOefNet217Ww+9+xMrW1aHB+6B78JCEisQ6Pd4vel2j+qhza2w/RvfRLf+iSDGpEx6dC0kImLh0wRwiNYNpOUht1Z6VM8unkoQDRrsnViMWubBAwrx85V3pPzqCpamouaICihmQmAxii3ebteN0zMzEzsgw/Bh+DZERMRI7EL5AHMVKuKvbIHJ87HdbPKgBb+8t/+27/8d//un3h4jjjiiCOOOMSRgD7iiCOO+Npgf/mXP15ttyezup4Fb6xTBhcCMZFDdEPBusLQl4vQUiepTbF4VWZQtZx3221K0TRXwQNCksTs2Dlmdt4xVcHXohiTcj03L+sobVY1sD2B2AMBvOP5bDKb1N65LnYxZiDKImjRDEsbp9LPDBG992YgoqWos+jLDKynnwFEhZgq58rHyj56xRlz+cgh7+u9zzmX7ucp/wInwV8LvaiThmJRx+zYwHoHZ8J+BVVW4APxXNhJBCxL96LOBhuNOA7Y3r1iehR+9mOLB7soss9ixQu9o+JA+o2OGwADo4tFaHyPbbzndGHDHr8yeABUymT3UrFRyToIUcft9O8O4zIIZXFUOg8aaIDBqWPYe1mgDkTowDaOHGqvgLa9q0d/tXoO3mlCYmK3XM6F0xribnO7ulsB1s5Pw3QyZ0aGFGhze7tbryUaAfu6rmcnipQMmma326xjmyaLk+X52enpeRcode1mvb57/QpSzjmRc86HFDttt1cz+t67F292svnpdVTKosxchVBOTVUL/yxZjCh4X7ye3ZA1aWPrHBfH53IhqqoqwweAXHTU7IrVRnmdiVU1hFA4ICUlIu+8DAghMFPbdYUFKCbOKaUQKiiW0IOQE8yyiogMesMevcF0T5qxSi4E9NAb0vYDPY4fQH/fH4RWH/+EhDwGbU8fFCLbtKRbDkK8ZyVgsPQAwL2RfBntkRUaJPB9Ogb3xzC8Z1Cctc0IMTh8/uTyD7/3/PmjxdRrapuchMPk5OKcHW03291uBZrPzy4mJydZdLte73bNNIRts1Gk6XJxen7W7bavP/vw7asX7PCdZ9968PQdNNzcXF9//vkXLz6eTScPnz45f/BEsr7+9JNPP/2kjd3Zxfnjx8g//ARAvjKXGAB+5cX/GoGD88FvjtMbpaqHfCGhTTwv6/rp1ez9Z5ff/+CbV4vJoqKalEHROU8UHFfF1plJwVxd+SrElJDIV6EKtXeemEMVvHNqJllMBJAMHeJQVZOjqhIiIJtaztKXZ1CZlFXyoO9EI2bPmESy5KzJRAnQ2JloTllyBgDuHdxBJKcUVcSHgFRUokIE6p2IpBib3bZYJGPsXCGg1cyAyA0FEF5VUkoqfatPH4qQm6SY26bUNxVUU9Us2XvHzEVxbGbT2cTMmmZXVxUitl3r2BFxTqlMVm3bIGIVah88EaWY0fo2DJJz13XkmL133lLXxZRKjsgQCJ2Zdl2azXwIdT2ZppQsIlExNgnWp66LcxQRkaEBaG9oQohmKppzni8Wk/nUOS8iKhJ8IO+BqdQ7EXJWy2bGtJhfPX188fTxo7PlYnu3ebNa3e3aFGV8+livd4aDAP2dZZ/3M5KKdCI5JTALPpTkKNM+6z8WowAiMaiZ9rFoIjg+UO5vvNwf0PPSg0k54PCA6aUDVKYMNIWSGu9rxQ6z1b2Dlxpkw86gzbLrktecmbL3kyp49g4JnUNyCMCMSIBmOcciys4ibc4AUr43eZ9C8FUVgufSits7co56Q3mHohBAT8LsbUxbpXY3A86//UE54ogjjjjil+FIQB9xxBFHfG14+3TynR9++Nd/8b16Nj2de5gA5hZB0Uwlp7bJMcbYdV2bYpdTRDRQ0ZxEsko2leCcYzZRRiXG0oI+eCIiZDSEyXRS1bNdE7Ohqyd+tqBValOOIoqgvfNtURIhABBh5f3JydI5il2rBi746WwK6MxI1XxwiFi0yUSFosWyHi7C58JSFQpSzbIIIjpH/QKm19SAonZt297zJzQAIKKcJcaYYpQsX1nJ/HrYWwj0/+z9asVM0dCQEE0NiVARURGhCEhH30xELOTFHjCIicFwON+R8oW9lceXOGQYFGiFvoWej6MDBdmeyRteHBWiRVM9MMJmxbPx/kLcAAAUpOfH9wrmcsCGe1Vz//uFfj64XLY/iF6ufFjvvAdR2Qjel3CPRicE3F8SG9hzHA8GQJN1SbZNk2U6nU49XjDazc3t9atrYn/mrvykntoc2aVdyu0qtbvV7ZuLJ8/QhWp2ckLsNqvm5q7dbpBotpyHxVykrqeTZrvZvn0dt+tqcVrNFn4yabarzz78Gc3P3n9yltzs49e3X9yJMnnvQwgioqLEFEJwzsVCBxOVwK6qUOqU66rqPWWIStakLNeL2WtKqW3bqqrn80Vx3kg5TSaT8u7YZpOd886llFJOkMB555hFtdg613UtKqIaquDYeed7ypbQzJyqSAKw4jAAe9UxDtabqCXMmPZK+wEjAV3MvA/V8QaGQKCGhooDL4x4MGJa3FOgV+aPLtM2ZCAKB31PRF9kc/c5oj3jXNJXBDDuStVEcoxtjO1yUv3hd9/7k+9/I2DDwLHrgP10PvO1j5u3ubkzk1BN69kJaN7crXabDWPYbJsuw9nl1dnVlUj84sc//uSjv6uCe/bet568/4GJrV9+8fLjn79+9SpMpk/fe3958cCYd6v1hz//SdM0p4+e4tVs+fqnOEjIv4KRx/kFd8Qvxe8Gc/1LoWX2LTS0AYLNmJ6cn3zw/vMPvvH4+eOzk5ln7Sh3zpAAzKDy1bSuJ1VlpoaGzvkq+BCqqnLe15MaDbJI27aOCZ0vuktmVxSUIJxyEslg5kMIwZuogTGR51CSZqYqSVQyM5Pj9W6DhERTZiZkS7mJXWq7Dil4751PKUrOCZGJwCzGrtntuqYpDwAFcI6YiRmbpomxA4OS2XrbNSKCgAhsgCLmnAveO+9jF7fbbRysqEr2S02QEAFiV4TMkFOSnFWlnL6BlUztrqmZSfsEFUnOwsakatrnddkhkQsBEFWBmMvTIGVBpMl05kJgx8jkQw0IVVWHEFxwAJRSbtvWsQvBV1XVdp1LyTmuQhWqKksuTgxFfopEgEUKq+zQezZRUEPEUjREaMikYDG2IIlDhYCMCCoekVHbtCOgeQg/+PbT8+Xy6cOL/+P/+uv/+29+2l1vY1YAyGM09SnPkTD9HRdB70FEVVV57wmx5M6LCB0AxieyZEEidiVLYWRFUXDvAqqJmQhJ/41u6KbLCGQkIiZiqshcXNR7BbQBmCAzSC9bL3P+kIYuB2Bi0HR5vWvR6U7VAdTB1RVPajefTbx3SBiC98Exu0kViLC0CAYgK90RcjYVAE05pxTRjAiKmBtMvKNpXXViiQIv6sAOUCF0eIyRI4444oivG0cC+ogjjjjia8NuWr/9swnEjlOkpsnrN6ldp65BUxPRnEoRbkopS9FeafnmjQQGJllEsmPvnWf2RiiFDSRzVe1Dxc4BcRTpRDhMFsvzarHML29f3d5u2lbvsSJ7jpaYptOpY1YR59xkOl0qKhAAEZLzDABd1xPQI3LOvX9lr27rG7hlESh+BQMpVoTBxTNSRYvUtJBZhdrrug4AVquV3eud9mujMG0D5Y290nVYi/XLKkJCQ9MifyYkOyiuHm1D6MtK5UH4PAhFcRQpj6LygckbtcqHYtGDg+g/VUAjWzt+eBRLIwzEuI0dAb+EkR8fhhR7trsnxA9MEg5J6+HT49/llHBYLvbEt+49RGC8sPdsPHr988H2Duh6ONhYjuv19ubmdrVykwVPZzNAjTlv1s3rV5+3uTu7vFxMZvV8ImeZwW02q7dv3qy7dHr14OTsdHF6EhwFg9u3t9vVnSEignewWJyR4grfpJSapplVdT2Z5tjumtVU04NlhdXie88ur28+3kUoEu2c+zaDKSdmbtsOAbz3WQTMKHJ/LVFHgVihoUvGpeQnij20Si/NK/p9yeK8K7aopb8TxrgrK3VVyT3xLTmb9SSummbJu2ZXbpBRQl8uq0gGAGLtyYIhtspRFQkxmOVezvYVDhoOVMswZEFsCOj9H2PQDSYt98idryro9ymKg3gcQvDwfduHgaoh2KjtLwerKjlG0O6P/+gP/vWffPfb7z2YYRt3jVqeT+eL5cTiNjYbyTGEMF+csg93qxVqrpzb7LbNrj1/cDW/fJABX//sJz/6j/9hsZw/evz08uFDI2pXq48/+vnm5s3lxeWz979VnV5YktXLl6+++FwkPX7nyeLZe82ddPlvv0TE3Mc/gH0+AgwQyYEpmDrAmnFa+fceX33j6YNvPnv49Gp5OQuBlMDQoWf07LwLnhwD5pgADRlIUbpOYld67cZtqaoBUdulruNV10VE9N4zMwF2qm3bqOQQqrqusvepOHGAeu+JUNWKwFhE0DEy7bqWHUvquhhj7GLXaRZTZezp1Zxz8WdHQDPNktq26boOh7ydD8xMiJhSFFXHvjQtNWQxzUlc0Qo7ZufIOXaO1XxVITEiOOfx/2fvzZokSZL7Tj3MzN3jyqMy6+hrunsOYAAC4GIJUARCrlBk922fuZ+nPw/wtp+AQpEV2ReSu0KAwGCAmenu6eqqysozDnc3M1XdB3P3iOxuADOzQzQxCBXprsjIyAgPdzN3t5/+9a9DQYIVnwH2g8lPSjGlrCp1XXvvDSCLiORQBee4dDot5yVmz84Vv+aSBibmqqpKVQoiMRIimSmxc96XK6OoIiIzhRAGEbSZDzBbLAiHCyD5UBXXYO+cc5SzDmJyK1lsx4wEKUdTSUkYBtcVUxU1zZmJkMhMUA2VS0qCyYEBmLAKM5AHZPvg2WxWfTyr7OJ8+X/9p7/84s3D3SYCFguwcvE7OIMd6TMAAKiKmdZ1NWuauq5LuUzOw13ZiIDNAIiYmRIiALB3Kl/tVlguGuWwQ2lCaAoAxW8dCRVRREqjzuG6rjZ0OjZKZiajDXRJ9oy1XaVtZRf7JFVYzoKpA/UEZtr1PaIBgkiu6ioEz87VdRUqj4hMzITMzEhaBjABcbl2CpgaqJoyQWBy7LOJUlVVs0aC39xn35vwP/oxOcYxjnGMYzyKI4A+xjGOcYxvLd6eVcQzk06293G73t2+bNc3u90DmTHAJIJFRAdICKKqIqbZ+4qYI6IaZiTvK/QeC8lFAARuZlVT+xB2bbvdbjNg1dTLi/Ps6m3OX7x5+7Db6Tcs2kwNkHg5nwfvwZSIqlDpgtRKza4rFs9VFYuo0zlXoHNpP8jMpS7Ye2emOeeUs5kxF9NJEBHnHDtOKUkWUCteuqpSVkSItNttVW0A07+Csml0GxxoJyoAFc8IVQPQUVhcBMOobGhF/oxMZkCiOjkZ4yCRLhhhcKuY5MkwrOcGP8TDz4cD9DyIicsScK8XhpEEWkGZWATFRUVW9OCTicf4eTa+20iT9zvnQG49YkNAGyk37j8TDzfogPEfcO5BGr//UgU4F6fIsmds7Dw1PNCieD1Ao3usPmzVZObBJrtt2N7fbO7gzC/IvPPVk8tnLty2u1baXXtzN3sScNH42bLOKsBG603c7tY3lTe3WC3mC0ySYt5s1t329uHammZe1c3q7DI0i9dvXm/Xm3xzqyer+epsfnLWx35386pr8XuX9Y8WtL1q25hTjDnn0v2PCAGh7yMRV1UlKqZqBo7LgreU26dpTw3fjGj8+ppTbtuemMws59x1PTOpaulKiABZcrFwRSRTHdIXg/cLqkhpKbrd7UwVRyuYIaljWsj+IfvGsQT+0UEdNc9QzHZHaduYNtg7ocBAfh8P2kdzaJ+BeJRVmPCymYJZKcsetudgrB+M8UKbJ6Bd3DbGpEx5fzUVz/TDj9/5N//qh7//vXeXHh7e3sQuPbm8mC9C3L5drx+8c7PZ3HFg57ebtcY29n3XtpLl2fN35+dnGuXq5eef/fivnj99dv7k4uz8OXPV3lz/5Md/c3f3cLI6f/HBR/XqXFPut5ubt2/eXH158fTps48/Mj+LP/9iXfJeXw38e3/8+ov/SeKwb0pp/ZreFpHQGWQCa5jPmvDsZPaHP/jOR+9dni+q2ivFLaIymSNjsMrRvK5yKh38Int2nolRRHJptTeysOBDVVVtlpRSTJGJ66qaz+Zmtttuu64F0/l83lVVSW2mnFSlqetStRP7PqUkqsBkjgQsVEFSe3d3t9tsc0yVD1UIiJhTjikzExETkpqCGaClnLNkIhgTsaZGSACEzoXga+c9M/tqllLqu975EHyoqlDqXJzzlVqzWAEM1j0l9cXOOedKGhiJHHOfU85ZVIu+1QBURVSJ0DkuHHl8E8flb9UkZ/LTjwpmxUGDmU2BmNn71PWp7/u+d8VFyFFKKcYoOXvnZ7NZKVkQEYeIgKUPJBKSaamgkZzFhJSAiQmzacq9SPbeMxGMCTbJ2XnvvQdVAEPJOSUA4lCVSwmZECJbTt1DhfzeZXPyRz98dr6Mu3tnmuNDq9pbyYTCdDk+xhRZsqhUVZjNmvl8DgAiSjRk3Q2H2o4y0ohocJpynLM89t8op3coPmlQALQqALBzjl0WFudEtaQsS14VzahcalQkZx3KtAyBhsvAcHFAA+tSFNDFajlj9KBoWVLMKUbJKaWub6s+OO8RsZk3TVOzY4fExLUPnh0BOMfOuVAFKikOHdIhzrFncoiKGSl4H5rgCe8ps1bNJ5988sknn/xjHIxjHOMYxzjGN8URQB/jGMc4xrcWSbjXTVDdbR9id9XdXef2QXNfeQ9EOWcobgxEhgQIBsaOfRXqpvZVRcTEgXzl6oaIR38GVc0pxe12q+sHQmqq2i9XoVmayJevv/ybH//s00/fPDy0h4LckUehAdR1/f4H752dnYrK1dWbt/dbQ8fsihBmWo2UBfJ2uwWA0bIAnHOlLpi4SKZARFWkV2XHYND3fdM0oQq7XQtmnstlyHKWIrwSiX0fU0qqpXUSQfG//qXDABSswDsYpZqGioBoaHueK6V34ojzoJgeQtl4QCjuBHagGJ+cRvaQ9Ss/jTAOB7o4eCyOjftGIegI32y0PsCxMLx8ZQVFmZ4Gg70hSVnyjcx3D4unDRsA+wQfR1HssLmjIOrQcOORXnv8MiP8pr2KGUbNauGbZak6EGdEgv13GaxDhi1WKBXb4B2HwCZ583Dz4DpdLprFcnVyEppqfXu3vrlv7x92vvG+plBRqH2dLhYzfftl7Lb312Ip08lZqKrFammo7W69fbhLXTo548XpaVM39LCBbdu2OyI8OTs9OTvd3N++vXobcvrB85NPP7xYd68/e7vddJ2OB7QQUAA0k7Zts+RikVk4EBGISM654OAJARMNxirMrGo5R0IkZuc4xqgqIsrMjtnAVFRUCpDLOdPUIbPYWBQkzZhTNitWzoAIjkvDqDylo8qOp4LMcS9tR7TJIMamQ7zPSeB0oPfq6P1keQRzDvImAIA22jvvzTeGtwYqvzUrmGmcCbifddNbjnJnA2DmMtWKzLp4hhPzxdni3/7rP/iXP/zwclXl3Xp9e3dyetbUoW83dzdvUspPn71b13NEEhFJferbu5ubnPXs/Onq2YvYddev3rz98jUTv//+B/PlKYd6e7959fLz6zevT1Znz979YHZ63rb9/c117lvV/OTiybP33l8slte3D3dvr3a7rX2Vnh/st18ovn6y+u+Edn/9MSCoX3Rj7eD/X42D9zA0UVUHNnf83pOz77379PvvP3t21qy8cdxYhoiWLOfcS+5BzbGrfAUGaiaq3nt2JJINFBF8obPeSUqx6x7uLcaYUhKRqqoW8/nDw73knFJ07Nm5dL92bleyQX2KXd82deOcQ7OS3TMEImTnHJMhrLc7RJ7Pl25BlQ/eObHB+b30POhTRERm9t4BgiE4x4655FCBBlccRGRyVDryIaloyin42rFDgJSzqnrn2DliVoVi8TxkDumgvggAEdVMRJOID66cE8q+zVkIwTnuYwSAqqpjTDElLSrXqip9d6NIETIrmOYMxX0ZsGS2S8ZLymmNHHtXMWIEAlDLKkPqS3IWVTdQeEgqZurYVXXFxEAlcaluVqv6qW+qI0YAVY2AkqWNKaVkYEycB6MGKhLsrImYnfeisuv7h/VO1Elrf/w7H81CvZx/8Zc/e3u97QXA8NHp6pcZ47/JkVPOMc2aZjabLZfLruuIxLki+0Uda1umvGlp2uFckUo/AtBmJVsxmqqVJLMaERbDFe88IiqYDrVRimBooCKSIxJ943ExtGLB0afcpZwBlJiYPYVqtaw8I4KZigoiZEntbkdEZipiMcbU92RAAGjovPPehRDK5YscO+ed94xACEwIyOhJHnYpk/SRyMfzj6F79d//OBzjGMc4xjH+zjgC6GMc4xjH+NbCwJqeNVjOsd/tVBS5CqGp65qZRXJZ0gIzEhkRDI3+yCE6ptJpkNhnANVsakVcKULdrt9u1in2TT1bLB2kmGGXOnnz5dXLL16/vdm1fbZRZ3u4SmDCugqnJyeIeH9/f3d/v932rpqxCAAODdLNzMx575yLfQQA59jMALBsdoHRzOwcSxYRUTVmMrMYoxlIlq5tzSxxqQW2sScb55y2u91ms8mDNcHfxZ4Pt3riIPsnsVRyTkj2wNZ1wsBQiBgBDYKgQXW6x7ClZx/ZgQgZi3Lt4IOGj5tIwf7Hqa3hVKN6oIqGiRyPoLD8dtAXTwroR+rlfQdD02JjMILEUZA9McABSk7IsAh1B8S0R9WP9+OEHMfvNRLzvSfICJoPtscO4OX40gE947gVQ2vC0s5uVvFiPq+qkPrddp2ZwdcV0eLk9AmDy51s1+v1+h4c183MTFxw52cnSePtzU27bS2pJlmdnNRNg4Tk6P7uPu225ALXTZjP69lCYtyt71VSv9vS+UnlXB38Uu1sEf7l955dr/tNl9489AWlMpGBoREhGZiqESJyaaRVjggAYCmQNzWFye582pN7aTDCkNIozshWupuBIQITIe4NZxARicrhGdTvQIUOENOk/ydEdEXhWN7WwGCQ5O+HzjigD50wxnnxaGLgPn8wydLhMYA+GEADfrVJLn2oEJ5Gpu5TIOPvH1lA73MRh++PhViZqoqk5Sz83vc/+F/++Pfff3GG2rfbjSM6Pz2BlB+ubx/u16uTExcaZG+aRaJJ3K7vt+t1PTs5vXzuZqvXL19dvX4jou+9/+Hq7Amxa3e7t1dXr15+WVX18xcp4nivAAAgAElEQVTvnF1cZoObq9evX31ZVf784vzdi4tmvtjd399dvVnf3Wn+evvBr8ySXy3+SUk17Rse/b0vnUj9lNAczrjFBwkB0OysqV6cLn7w3tOPX1y8d7H01lm7jRJTyQmCiSY1QUB1VlzTmTkEX9zSDQIREGHwIXjvg4fSYzBlF4KIIKL3LvigY7bN+4qdh8KXmYgoS+5jVwzfEYGQGAmYyDvyrnhGZcmenWcXnHdMhFiUngXVmVkB0ETk2JEjYmLHU62KmpVMVZnehmCAXOoY1IKvSnvSmKJkKdbw7BhxECyrCeK+tMJUy0tETFSdCjviyabcLMaEaM5xyT6FUKlaueYSATMbgIqJKDAylVIUBTUsGuokaEWijqWORbISE6KBZDGLIJoHEyHJWSSn8QoWU+nuSKWDKSAWGyEAFRFJOasQYRWqIlBPOYnoyNmBmFLKqkZEo1VI+U4gIF3XbzZbRG8YnoTwvWczzE8Y4adf3r+82USAXByg8VGOeRyHcPD4V8te/yPHr+cTd9vtw/190zQI4ByL5L6PZoZIBmhjxhlLDwMRMyNEyRkOblEAhivSwX0NDFVPJUtaXP8RiUjH5HYx2MEp8zkkKQkABzO0gy9rYLs+32+7u80ue46MjWeEyjF7R9575xgRRHPwzgYtgmVUNkEVUwM10JyTmki5saByx8m+aLERjZynELGXjhuUiExw9/8grX4tu/oYxzjGMY7xq8URQB/jGMc4xrcTf/qnf5pgxwtbzhoz6Q3qelmH0DSLUFfOe0LwlXOVR2ZwDESldh1UZP2gXWugCKCp267XfYyiulqtvPcq0m8f2vVd33a0lNq5zf2dcYXV6ur1m+u3d7vuK5hlWrCZc1wFV4Ww3W5evX693e2ymB8LMMuisiibiJmIdOgx6Ia1tyoAqKokdWPLNTUjojhZFYjFLhaD6CL4Kr8hYkRQ1e1ut91uUx5+9U1rM/xmJDQC1ZHroRX3BxpoX/lDZDpApEjFlpImBo24t73YU2gYFG1cVstF82tTh7/DtdrIayf6PC2DDylzYYB4+EnDvtgrmoeOiFPzwEGvjDis2HWCgY8sFBDoQIpd3kFH1+29phlgLJ7d70HDUQw/sej95g37ctiNI14u5fDTrhgBKD4iAiMoV1BTnVXczJez5bKqgb3kFLebNXFYUZjNV0+eE/pwd3sdr7sQ6qqqZrMZeT4/v2QM97d33XaT+iszXa5O6tkcfRXNbe9u7+9vFeEyvH95cVEzzeu6262vXn4OuQNkEXUOtX/47rPZ9Xcv122Oer/Ng5y/uGToOEixKBydLzYyquac896rammSWbo8lXp5QDRVY/Oep90VQgCAYmheDmV5vtTuO3BEVLJIqipFn4gIAE4ZAIhpAPem5aOLMppH8aMrjcYG+wsiZhtEa2PSobCGKcswwgWiSXM9zC8dyx8OyfHBCEJEtKKmH9jCo1mII3MAAtO9MH4/qoYJMQ6ecfyNY8XU1HL67rsX/+u/+aMffvTOopb+4R4Rv/OdDwO7m7dv+106WV48f/F+AuxSBu01bbcPN7fXb2ez1dP3PmjOn2ofb67eqsrFs2fP3n2R+q5b397dvL27vZ/NZh9++PHy5Axy7jYPd9evt9uHxdm7q+dP69Mz2WzfvPx8fX1HqlUI33Bi+UVjj1/H+CfFnUt8Rbn+DwaOp2g7zH1pOQkpKAEwgAN472zxu995/lsfvnNSM6eHfntvqUPNJQHIzvnK+6qqqqqu66ZpQgjlMRN575umYS6ck6bJWBzYS61MVYWcc4yxamofauIgaoDkg0cCJKxqX5AZESIjEFlSUyPnSnO8zXqdUwKAuqqCD0xsKqbZABBpdIUCwMESV0SLGhuwMFdRURMBSOxL2RCmnLMkKJgaHTmHhGTmmLCwMwAV9d6xd+x9ztHMgvciklJquz4ErHwjGgsGNkBDcMjlilzSXGhQh1DO08EzqI8pFZ+MFOPQhq5YKjCVw+W9F8mxizDkhwhK37kUNYOBxq4rfR0kqkgxpAIwSbFPKZXeqqqWUo5dLzmXWW0gOaUYY99HU3Xez2fz9cP9brsFBMfeeQdlQzy3bWdmdV2VS+FiMUsp7bY7BcMhNdyrWtfnU1f93ndOnz+Z/ee/8u1/3mwEWoU4nuNKV97DQTn+/+tT8heaAP+48Wv7xIeHByRaLBYGpiqbzWa73akKki+kHkzMDNmVVquWk5UWBMwIpdEfAKKplFuYr27oN2QpS+LBYHDhgODZOx59mWi8wXjU/UINdl2+uW9fXt3MCRqEReUWdZg3VVNX81k9n9d1FRoX5ideLZtlBEOYkZUUvUnWlFIu96NZRSyr9m0U6UxKB+xsROQDVw/+7GJW8dqEW1W8/XXt7WMc4xjHOMavEEcAfYxjHOMY306cNOllO/v+Yntx8cRDzo04JseOyaOpqYrKpu1ksymARiR3bas5O0JLiUFDcIRIaADofWCzru37rifiup7VVSMiznnnPLqK6qVfXISXW4CiMir/s4IJp1VFqKqqqYEwpdS1nYhKtj72kjIYMJOKGEAIQVRzzkXhGWMUVUIMIUwC3tI0raxMymIVihZUFQFE1QCYi3ypmBgQAOaiQEvZRCdk9qsFMSMSIsHoVVB+3NttTGRwpM8Hdc808LIR4A3PFmORkgyArwFoOFD9HqihAQah1gSaoXQRHGjGAZkGNDrgwftPHwWF5SOKDHt86dcErjCSvv0fEREY62S5a6MHB0yv2XtPDx3qYBRFDwSRDuXPiAOrnhh32YBCnnHUex9uNCAwkBGllA1weXr+3vOLzZtP79dr2u522zZ2/erktJnPL0KFzl9ffXl3/2a1XFSVTymL2un5RfD17durFPu+7di5uXP1bLbIkvt+t9msH9bkXs8XC0B0VeDsFeH2/u7k9Ekzm0HfXt2+ffeDs3/92+8l8Zv42ef3gkzO+dExRgp67roOAJqmKZXHYMjM7DinXJB0VVXOcVEEi0qMQymA9x7AYowFaheWjcUCVUREnCtWM4PxNLMrLcCm1yAioGnZsQYiwkTOOdGhpL0UIhCRjQC6DKyhgr4IzEa7lUdqwAOFcsEO45D9BnozdrnEaYDQ12fjNPLG84mhmaoBjahiTFyMGYzxU20c2AaAqHZ+vvoXv/XhH/3BD+Y1b+9v2Ozk9KxazG+/fNV3sWkWs/mq66RZLfq+7du+366vr942s/nFs2erk5N+s/nRX/23h4e7F0+fPHv2tOS92r7d7NbO0/d/8DvVfKmSr9++vn57Vdf1hx99dHp5UbPfvH7z8m//NvexqeerFYdwdVjfcIxfPspoKlpLCwAO4HRWffDs9LvvPPnw2enCa4UanPrTBcEMTIkde++rylXeBRd8KOGcKw+YqcwsVRXJSCQImhMRseemqbxziNT3HXNYNA0QITEwe/bIjIQARoTofHEujilqVmIiKA0MuukEVwpxEFFMi/VEKU0Qs5TjcMKj0g5YASCmBADMbKZauo+Oc5lZzSxLFpFo5tgF73fbrCLTeXMwoAEIPjAzAuYcTTUW1w7V2LWx61LfT4ULKScwrUIFYJolpYgG7AgQVLSPfTntppwRiJhVBIptFCCAqUnpMKgqOcUUY/FhAIA+9lmSH2wQZChvYpeipJhTSkRQUgBmKqoqOuSU0+BbjYgGlpICcFM3ooqAKQmRq+oZIs0X88V8Xm4YDCGEpkBP0YwIzldqQM4F7xHRJIMKMc2bWsllcsuTpQvN8mT115+/+tnr+y9vooxZ6oPbmCk/dijP/2cRIiKSiZCdr+ua2RVAjEQDcZYxi4iAiEYEJQtOhICoOtyEHPitTVGuPl/9SMRpLIMhIpScxGF2/CtRjlRSSIbGznkKqJpTu0sa27jz3dZv7r1zWNd+sZw7R8xAjG7cxlJTEKgKVV3yL2CoUyGW2niiAGBGR2616n29uVlrK9bkTz75d5988h9+zbv+GMc4xjGO8YvFEUAf4xjHOMa3Ex7yd84zA8zr4BVsPgMsqqokKebYxxi7vo+xN8mSc86p3bVgFkIono+qFTtm5qquHDMAdF2nZkiuqqrgAzKBmap5YG5O3PK8l7/dtv3hwmDCkMUioK6r2Xxe1fV2uxVR74OATrJWInKESFTXTYwxxr60FjQAS2kiTQBIIzxmZjMzERpXQThqMYnZOV+gGwCEEBBJVQAOepT9aovHQZg5cF2YUCjio65+MMoxJ0q2F/CO5Az2y7WJ1BWrhPF72N6eYjBjOFikFWsSHD6IxnWdjfy6EMFJUFwWf+PfTd/l8X4dJMqjyvlx6fEjm+lpX48vIAQbOgnquE4/3Nr9Hh8J9cHemPbDwWttYugABVrCaPox1vuO7zhszLBUVVNkrlYnpO32jrrtevdwi6lF6RZnT7lZnV4+N6T1wx2BrLebXdtVYbaYu3o2Ozm/6NvdZn2zXT+IapglRJqtTjjUOcZ+t7bchWZez+aL1erk/OzNm1frtl0QVVU9b+Zptz118+9ezn/67OTt9hp8IOcKCSrtuZhdkfk754avUlIXiEUIyc5VVXDOle9fzDQRwTkOoQIwHmMaaUWqKSLeB0QS0WHklBlhVmSVOWVmAkQp9eUAqkMtNAOX4zKaq5KRok6HA8hQAcBKOTUeHPdxZBweoPLxB2Nm/9r99BnksGr7HAx85V0n5f4o6jcYDKMPPnli0KUcYajZRhumVOXd9z989w9+6+OLZbO+u7HUny7rqq7XDw8x5Wa+dK4CdKBMxqyQd127bheLk+XZ5eL0POd4c/Mmt+vVarE8PanqkNrNZnu33W6q2eLk5KxZLGOK97dXNzdXMeWzi2erp89q7x6u337+05/s7u5OTs+bkydz6V31czvcccf4B2N/hplkp0OzMQdWIZzP63cvV7/1nct3L1ZPlnVNVpFWjLO69t4hIrvAIbhQFTuLqgrBF/cLLq3SnCPi0UOAGJkNTFQIEYiLfpOwSJvJVyGLAiKWen4iNS0TzcxEVDX3facqzjEhg2HOCRCL/Q4TEbDkXCxvxzxkURvLlAiUlEvSSMrLhtNi8Zgy5xxozkjlfcpoFyRhjn0UEQQqaSBELDUDOQQmAkRJUVVKKtTUur5T1XaDrniIALZdm1MKIRCimeaYAIb0rUju+77kUlNO5cRVWvuWxJWIiKaCAIdWcTFNPr997LNm58hMRHPOwsTBVzmrZMk5EaJjcuWiryZSukEiGBCSY1c8pp0hEnrnZEjfQeVcZcbMi+VysZh3bZdyFlNmBoPSGRIJmrrmGIy4mc2IUGK0HAmhCrUiZqTTMF+enj198fT5i7OTv/6i//PPHtrUZ5tg8zgKJxn/12XRv8mhpiKiprV3s/m8qqsqJjXgIQ0DxQJlzLejsjOwclcEACpaLgYlufL1jOPfq4BWMKMh91yaSJsO+dRHx8EABCAaREAgbmbVyiN2LWomE5OUuiyxA9SudTknH5z35L13zMwICoBAREyOyRERIQ99P6fiNQMzYwYkBFJervow//R+J5jpstvtjvTjGMc4xjG+tTiego9xjGMc49uJhjprTQOn9YPJFuK67zZ93/bdTkVyjH3XETEApj5KFjNg50NVN1VFjtk75wP74ELlq4qZEYmbPLk6KJH3nogRGZAhzNXNXr29e/nqjYkerAhw4IYIxDCb1Ser5enJabtrfVWdnp+1UbKYI0YwUSkd1rwPMcbYh0LZiDmlJDkP+k0Ak2Gt4pjNLKVUXoYAOecsAswh+LoOMaacs/da11VZFu3aFhGNENSgrG9/qaUjYkFgJgpqQHvpMZIpOySj0ioPABAUFY0IDQyVFBWLIW8puN4TN4GRXQMXF4NpD5b3xhFKjzFKUA2AJig8vhRHIaoB4LRyggkPjha94yEaPmakwgP2/fpycBQuT6vvR0/AV/5kIsgDI//ajn5k7QH7zRvpsw4CpCGHMQmoR2Utwoij9m0uEdAsZYlJjN3s9Mw7ar3v1nep295evVJ0S99U9Wx1dlHVzXZ9t9vem7SVTwTcNPPZYulD2G5v+76LObu+r2erUM/qZhHb3ebu7W6zzgp1M1+sVgbLXYq319dt14eqWq1ONg8P3suT2n10Mf/Ry5u7PrYxdn2fUqqbZjKWQcSi3C+HV0RFJPgAOAjNAFBFRvcWNNMY+xgjDahLpmFwuG7PSRCJGAdeq0bjYFPTLFmNplaHalpMA1R0yjiISBFWj57sMLzgsdHmqHKekhrjMLDDF0wH+SBrgY9SP7YfhCNhPMjdHAylccgQ4sGfT6mQEUGXpwxsaEiFqu++8+wPfvjdH3z4gqXr2t3Jsm6amZmlmOrZwrsgGbJA04TUtu16LX2qQjM/WczOLrPo3c317dWb1SzMlqv5cm4I7W5zc/WGfXV6fnFydpZVrq7e3N9dA8D508vV5dNmtli/vXr76nXcdauTs9Mnl7Q8o+29fEPG6zefW/3/jQPzDQBAQAIs9HlJ8Nvfufz+B09fnC9mHmrKlcPgKDji4HxVhapmXwE7NUySTSVUROzYBTCLWWJsnSNmUlEffFXVRAwAhOCcN4P1euuodezU1DGkvlczDqHybCAm2USJmdFS20lOOcecE4Kpc9mgTCEiAuLCmDORZMmaVaWcZVWkVAuFKgBAyjF1UUpWFREMYh8JwTsPxR3efO7a4qGBCMTsnRPRXd8VUOvY79q273rnHICpmXiHRGCQUm+qTJxTyjmVjnwxJlN1xFVVtbtd13WlZoiZUk4I6LxDGDoGmFnOuZj/OOfrpgbEwYRZBMBEFBGWyxUiAWLX90W1TYQE1Ld9n/qUIhH6UBH5Yo8yY0IDAEW1Yv5DzgFAIYCeXVXXACBmSaUgwqEZY+muwBRC8M4TU+WDV1GzqqqQymkWiJAcp5SalFbLpWOWlDT2KhkNRC0ZGPtVmL33weJ3/8Xvfuejn9zc/Z9/8/P11UM6GHvTQJwY9GH8ps9lM9UcY79YLldNc7I6QeQJQNvgpWbl6CCRigAg8WA4Xu7fsCgAfjEAbThYRU1NCEuXwRhd33dduwMAsEMDDgQAQesMegAFPVnN3z2d+9RDipIjFPWy5FJqdHNzCwDMXNe1846YnHdFeOFZmZWZGQcDKy6uVgjeu1lde1eaghrOZ75aNCHcb/rr62bhFI5xjGMc4xjfUhwB9DGOcYxjfDthqTcEphB3D5vN2357F/t1Tp1K5lIOaQZqhFj5gAERiV0IVd3M5sAETIjsQuVCoKHBkY50yUQkG6iIGmaBrIAhYW0/+enPPv3s8yRisCdRRTGEAKA2n80Wi4WaJZEs6pyr0HsDR2SmOWfnAztXLHERoYjUmNk7VzSeBYVLkiLvLda0E8gz1aqqiuzLOQ7BeZ/NzDkGwJQTtK2pWukz86vFyIYNFAxBi8ySbEClgoqGqKPAGbBo59SMyAgRB21dKTgt/XYGMfUgjjQaZJyD6pkQEW347wDJWekLhUSGVkThxeh3EI2qDjJkIyIFHNrRAZSF4uiSMfWrO4DJh0Rx4tTj6nv43ENYbKMv8PQ3w3sYTlrZAwE24oG79P4rHaJL2xP2aac/Nv/9Grse9bAGkvqu3+12MeUm+PrkrKnqNoT19evtdoO3bznUzdIck1+dGGjMMff9drupna+891Xjgqtmc9lZSjFuN6qwDI1rKgTouyam1LVd1+6avjHC2WzZbnaSUtf289X85vo6p7SoTn74wdmPX9/9l5+83W1TFFPTsvWmWhycc86qCoAhVCKSUvbOIaKaIhKYZcnMxQbWqUrOqWg2B7tYGwE9DtLjklMoOKZA/wKJB1cYg1K5jFj6eUrRVhtYafZV2K+oqhoi2ui3XISGj8y8y3iYch64n+y4l7EPuY5piI1s+PBg79Msozh/evdBbA97BTSMYu6BW09MHBHRBh31XgGtSgiVg9//7Y//px9+/OJs0a/f1IFXyyWhtm1HLsyaRexiFmFkJlrfvd2u79nR6uyyWsw4NDdvXl1fXWnqXzy7rGYL513b7m5v79pd984Hz8+fXCLC7dWbN2/eINPls+fP33mPQtXe3n35+ae7h/uLy4vL5y+q2fI+att2u+3uMWTBxw9+1ZPSP6V4VDTxywaCIhihzT2/c7r4+NmTD985fXY6n3kMbExDwXwZ9EBkSGJgamJa2vqZQcoCEKmkAGHIQoZQFQ+oDOCc865S0ZxTTtlXVXB+SOhkIecY0eRAfSwpqaS+S6lPOVXeM3Pxhsp5tFZnFi3tPanvupSjmHrvHTszzcXgWTIipJhEREVMzVTLBESEjP3BDDIR7Qtx9o6IRKTvYxVCSQy3u7brOyLKKfUxVqFyzhOTiIBZqRxCBOc9GOSUEDArIPSiCoOnf07JRLRchInQsDRN3SNGdq50UAQiX1UeABByygbYLJYIiH3fLJaIqAY0lM9YzilLDiGwc0RsZkQcvC+OIZ65fIpkKYJbRnLOhapSs6xiWJyuSIpdQsnQMfnSxBWGqwSWSyMMvkNF7y4qOeeqrghAUrJUmUixKVFA8hU4b+QjuI/evfzf/7d/+5/+4qd//uOXn726a2P+eyfnbzp6HsJUtO86Uw2hapq6jzGmkiUt2WsojYiHiw4w4NAhsyQ7B/lC6fPxeKc96io7PTk1gTTF4eqZJU83JTYlLMfAqW9xFtns+j6KGTjHVWg8zwZXGtWsIlrG19CbAdAQsHS1RswREw0VNXujp2I1woSeuTQzJAactzLr+rZVy0/6Ksd/DqfxYxzjGMf4HzSOAPoYxzjGMb6dMI0IFNDF7mG7ud083OW0AxNG5FA5HyhUpYS2CoHZETsm9qGq60ZAxcwMXClJlKSDIaMU7KOiZqaEbUzbNm77jG7uZpvPfvbZl69e59F9YSINAwkDmM9n8/ms7brNdrdr20wOwCFyWduLiHNmajH2pjYqdk1EJu7mnCNiNCgvICIb1wammlW99977LEKljpKZCEMIIpJzkpwly0hmf0kUcvhyM9hT2MHdYjADIQJEIBxMDQ20dN8xMDMqrRQRFRWp2HRaqfk01BHg2h5Aj9x58PqFSZmMAAOhVkWkgttQEalYowx95Q0RSUmJSHFyxhjErcMbPQLQozB6r5T+KoCGqZXgyImt4Emb9g3sQaSN2BlHifIATMt7lfTGo928f2sAGJs0Yukl91XnR3v0YACfLKltd+v7+7Q7U3Jc1W7ZkAsx9kbUru9T3509fdGcXDbL0ydPn89PVvc3V9eff8oojEmS7Xb92ZPLerbYbh7a3ebh/pbDLGUl5ubkCfu63Ty0m4ecOgEk509X5+uHu9u7O/YeEFKMp0v47acXrx+6n7+5vnnoc0Jkjn00MBrbP/Z9H2Myg9nMVC2llGIsDKWMFlHhYaHrSt1CYcfe+xEOl7E2aNsLzj4IGpMg+6MsKgbmnCtqNaJRrF9scBBFzWw/+0pjT52aV06TehgzZVSWY7b/7P0xGQFxkelPw8MOxtgEmqdfHKZFYGiquR8c+1TJmIQYNdYwAutiHaKN5w9eXP7x//zD771/WaVNn9Pl8yeS+rv1Oqe0Wi7bmPo+N/VsXjebu+vdw21VOT9fqK+Fa+26zc2Npfji2fOzi0s0WN8/3Fy92W3699//+PT5eyG4+zevfvbXPwrz+dP3Pjp/5z2qq/b1lz/6y//abzYnJydnTy/np0/Ahe3Ny7dffnF/c12aah7syK88+A2GF/Yr0Wc8IExGYExQO7xYNd95fv67331vWWHDBpINzQBEISMTU1bFLGIRSI3IALxzhC72SVJOjrz3hGSiKirmqopMNOZERN55qKqub1OKqgo+EKJqAcrJBVWVnNLolo6Sc06x73Y5JdWMs7l5Z2opp5SzmRETkyu8GhHbbpdSVLC6rqtQA0LKOeUsKQNAabhnBjknyWKqzjECZh3cn3POpQyia3skdNkjljIFcc6hqIkkzWIqon2KbdepgVcotvKIUHw8vPccKsjZVcrEJekV2LtgIpIlS84U0LHzwRePjiGBKhlz8s5XIWTJAMDes3PltJZSVoPF6gQAXeybZua9K/UWiBB8QfkQ6gpLxVLOCBBCMFUEaOqGmABUUs4pxz4hIRN777JIUiHHpUfxcAlDGxot4KC0BRyg9FA4ZcZMQ1tjFZE8ZK6QgNhEwMCAgNiHSgz6lDW1T5azf/cn/2qxWNQhqPzs1fXDtov6zfMTf/lR/U8zDERkt2tjSqVzACKl1BEhElm5RqsaACGSjIZgxe+l9IJGBEQ1g+KGNsRw3vsGWQDaaMFR6tVAsuSUZLy3efwOOPwFIILlrA/b7n7TrpuAzsIshKoenXfGjhSmopaytN1ORQwGjxFVHdzEhrYWeziOAKaqkouhFjFRs9PZrl23Jtpgnd0/j8FwjGMc4xj/Q8YRQB/jGMc4xrcQ9skn/3Xdr+eQldVSNaucPzc7QwA2InbeVb6eixoAVHVdFpauLDEBrW81RQSRfpd3ySQVBJVSUlNELPfwQNg9bG6ub6/ut9GC+dXd7Z3pACqtKCRHz76CmJaLRV03N7d3r16/+fL1G3CVIZshgqnkPsaCwg2MiJi4YLKUExcXTlViQsAcc1mr+BCKmIuITLXrOuccO6ciRT0jImXJXdeNmW0225QzEplqAV9/Ryebw3gk5yzOuoWojQpQKqzPALXgMUIiHgEdTcAOAArWJ0JChLEF3944ulDnkbROUPiQ6o0bhTDZQ48bV8gmEZnpXi180A6uAOgCIIpXc/l2hUJOfHCEzpOs1gYGPMrvBpMDG9doEy4eZbOw59oAI9QufzG+cHK1/sqXs0OdLE4K8ML3VccvdSCg3aupB5bqIecUd5v7qy9+Vj898adP2DfI4fn7313fvb19+2q7Xl+/+fLdZt7vOMwX9Wxmdmbtpttud69fMvuqns/CsmYyBDW7udvc391ePK0WqyUSBcdosl3fb9ttaOoni271xQgAACAASURBVKdN1ZhojGm9fgiV7yTm1K0o/8nvffzp67uH7tPPrltlZmMiLCMWAKqqYmZVYybH5L3HQdesg4Z86EtJNoqAh3KEMbtAzKaaB0+P4q0xIKoxvzC4spgZITGzqqhp3/dl/Rxjj0TOexEpK/xSOK9FrgkAClbG48ABxm0DnMDxIw5cBMgHiYID9/JxgI1HsDwcAHoZ/o//rPxzKI3fT8lxyIw67PE3aGUaOcLlSfMnf/jDD888trc59ecny6YKDw9tVYXlYuHYX1/fn52eLZomde26vXcVg2NDIvIq9vOf/TS127Ozs/Onlwjw8uefvf7yFaq9++67J2dPoNvdvnm4u76uq+bddz5YPHlKQHev3/zkL/48tdvT87OLi8t6NsPK3715++Vnn968vWKmR7P4GP9QjD1eh5MIg60q93RV/+C9Fy9O59ptul6FjcmYwTEE5uBdjDnGTMSmRs4TsyKoCCjM57MQvHOEMDaNJSTm9QMXE2PvPQCIauw7RFjM5tKn3WabYsySRXKShERVHQYhJyKYqUrsO0IMwXebreQcY/QhOO/Gzp+Yswwpo0FzaantWh8QCYiAcP2wEckIGKqAzDklg2JHy1Rqf4gA0as67wmx6pOZImIIlXOuZGgBIOY02+caTc0ce0Q6vHyxc0ycUjKwBXEIAQFTTDT2DEwp5pzreoaIKaVi9+y9zznFFHNOTTNbLhYxRkT0IZQ2dCJZ1VRhuAoyGwARusAppywJDb333gfJWUX92E7YEasJArimATPJ2XlgNT9THYpsVCWDMjoeXIaZD65+Y9IVLeXMZIE5ptzHaKZ13TjHKpJyTimVtIFnlw2yaEqC6ICpzVHVVESRHUKF6fd/+6OL8/OnT5783//lR//vf/tZb5ABHjss/LOhzwCAmEVvbu9Ozs5PT89iTO1ud397izh0vN3fPJQbP+LhFmuszYHxSgCqKlrqwIh5vNUYaS+MCW+iYfeaDpcMFdBcBjO5oKqgeng9GHPdkEQ3u/j66s7H/iTg6bw6Xcxms2pWV3XlAY0ImJHJiLFpFqUwkAFMTXIGKNOEVU1Ey+DSYRhK38exDAfEVGIbLGdDaZji0YLjGMc4xjG+tTgC6GMc4xjH+BbiLy4vf++nV//xd9hUkWC2WLDzltXEUIHJswsuVAqgBoYFMWnOAhoti6ReczTJqAk0m6RCnXa7XUzRVKtQ1U3dzGZN8KvFAl19ve5f3ty2bRycaREH4060shggACaoq8p7v9nuNttd10VXOUMTURyqIsUMUA0JRTRBxr4/8AcYUCkCTABazRCxWNaaasoZi0lukUERwABVtVgQ7na7lOLBrvqFJYcDMcWhkBipLJ1w9DcoRgOjYy8Vpj/8esRjZeVPdCj4HEHbQGoBwAbnXRvsBmzy6IDhJXj4wGD0HAAcAfQBFJykyiM9BKDB63mvJzUVGGn3qGW2ATIPbrqHm/po9xVGPDKA/Q4dt2Hw8JjsHAqf3u+Pyfp6VMweQHcwACKD4egbjl26yu6YRNrj8ZkANFSVrwOl9m5z3bKm+cllPT/xoQoKbtdiFyXnLz//6eL0/OTpswpXkrNvZrGPuW1Ve0Ok7YZ95apmtsTTXvq+2zzcMup8sTIVHyryIXa7uHlYLlfeVy5UddO07cNs1nimGOX1q5fz0+e/9d6Tl7e7Tq7vWoMRJZVGf0XEp2o4tm0CABnakWHhxRNrdszeO2ZXBlQRkDnnp/Zlo88GqlnOeRz5w+ARFQRkZjVS1dKIjJBk2oc6Ss9Ry8yCEfUXI4CRXBUsTAeu48MB2Q8qG04pBx7gSDhYRU/keZp4enA0x+cPxdaHAPrw370aek+fwcpgJbTlcvb+87Pf+fhyzp0D5xwQ6G67ibF3IQDRw3bXzBf1fJ4k7rr70LDnkJMAOUd0+/YqdrvVcv7k8gk4fvPq5etXL0Hl7PzJ6nQJlvrtZnt/Jzk9ff7O8vTUMzzcvHn7xReW8nJxcn75dHVx4UMVH25ff/q3cbdezJpZ03wlkXSMvzdwfyIBY7Ta4fm8enG2OKnJaR83kTyBI2EgBmFCP4jgRaQkY6qqciEgoWYRkXYHkn3wDgDKFCMqydeqeM2klFSkj5EIvHOq0vd9zklEVbKYiCq7wpBNVdSACRmRB9xmKiKmxMSOmalkbYnYOWcGJeFUev4hMRIhMbFD5rqJ5WLH3gFizhkQiCn4wFRcsRgAVdW5YrthpoYIPvhiXV1k4BXAkKnNGaBwYIdIACaqBoO3FQCklACg9F1ApFy4GyGzE8k5Ze8rACgmVwCACN6sNjPT4H0VKldlA2MuX4QAQEVFVNXKM2oKYMaAyOyQgZkdEKMBgpiAFT961dItMKowMwEyERbLlSEdOrh4mNlgE6RaknFDDtMsS04pi2QhKhRbc04pohmIIKHklGM0MyZijyoliVAksyAipoZgtWdgrgBWs8XZYjmv6tp7BvyrT1/fbHYwpWcfDdTf4NqFIRCL7r6LfW9mpTRHTUvycDKCUtVyx1haeOqIpPdTGQDNQBUQwFD2aWWb6h0KtUZmKNf8vQWHohVRdbGGK1n0Rwns8o+ItW1uu7QNDH2W2HVdW1d+VodZUwXPPjjvyDnyjth558gzu2GE+ZI2JeYhWTQW4phZ8csqKX40SOQTVxj0epfaTmZAf/rv//3/8Wd/9o95aI5xjGMc4xgljgD6GMc4xjG+hdjN7c8uf+eF/RgAHfv5Yl4vlnnXap81q/ceySkAI4nprt3FlEoNcU69pMQIZCopeUbPoCrl1n/X97tdm2JczOfo/MJVJ2fL1fkz8M1Pfn712du/TNmSDPjQDogUAjBhYKyDd8x9jFmUiEPwagiaCQGZg/dFNgVEWWQozkUsixwb+h8WWIuAA4xW1RjjoTPDQPcQjDGEqiiCY4xd17XtLsY0iUN/0ZhUuog2yJ2pWF9yMdtFBFViInZl1X0Ip0fnw73WFw8FvLCHxOWpSUQMI42GibHCaI8x0kKYNKcTgGYalbPDqqws71XE9iWxA3De+zAOque9UhXHZb8ZjmYdoyQVBj30aHJCNqw8h4U5juvJPftWVTWZkPYIGgmwSBH30iewvSga4WDn7fs9AhyuOG38bdHcW4DcNE0zaxgepNvs7oqk3gMF36zmp09VtNveb9cPBkKeREUBm+Wq+Lrkvo8p6mbTzMBXTWgWF8/81asvdus7TS2BGLlQ1YvVSba83dx3fReqOTkXQr2+f4vWLObLjbW3dxuz6+9cLn/vo2frTv7q5X3CQETsuIAe59xATnTIXZhZ6Y/EzI6d8y7nnFIipOJT6pwHgJylYBfnWAeL2BFsGpYF88CXRcouEpGihS/yelUZ3SqcmYHquFNxSBLsx+DQSA0BiYogfUoajMLmgr7Hg6sqogBFHz9K5qeDNmji9sxgRNjTsS/njDEFs//VOGEm0/EhO4IjnxqkdwZg7PDFxckf/vDj56e+dtkhoKFmy2LFl6Tv4263e/edCwDtunWfd95THzO7yoUAmjf3N7Pan56f+io83N6+fPlF33eXTy8vnj8lhu39/W69Vs2Lk8XZ5SUxtQ83t19+eX/1Zr48e/Ls2cmTU1dVfdfd/fzz7f3NvJlfPq1ns5vxOB1iaHv8429k/Ap4btIyApgRmCdb1e5y1Tw9WXDuUsymqZo36AKMpwrg4v6MSQQKqGL0nh07dSqqlsVEYJx65TRJTM2sAYOYkopkMOdpPp8HH8wUDUoGSBlBsfE+hKqqqixJJKuI9847l3Mq7sYAroiFmR0CxFRsPVxVNQCQcnbOBe/rutaS6UFCZmJHRIgEhMXyqrjlEJJzjhBBrQicswgNmc1SZ4NMJCp9SlkSENZV5bwHxHa3K/cAzjliQvr/2HuzbUuS40rMzHyKiDPd+WbWBLIwNAhQ3U2ySa2ltaSlr2n9Bn+j+xP6B9SPrQc96EHTUktqtgAQBRQqMyvvdMaIcHcz04NHnHvuzaxCAcTAYp+9VmVlnpg93CPCt23bRjFGUfXOF6Iw1KEMW2MdGVNhHVMU0VB5Vc+ZmQUUg7eEyMxd3zvnvPPWkjDnlBVVVWOKxhhjrPEBNAOzNSSqOUUkFOXY94BqrPHBKXPse0QUEc4x9X3OkTl3fZ9Tss7VVair2hAVUnh461OJjimLCpdqd8Upmg0Za8kSpZRi34sqIeY+EgDkHHct9zH7zvvAwjn2qiJkgJmziIw2UCKQGQEMUWWNdZZV0eKsri5OvjcJofZuvftfdm3Xs+T3ENC/XSf/NqE87nNO5bXSNE0zmVgfhuCnGbJzhtoGCsaaQkAPD/XxC6eU4SVrsVjKpFzeJUWZjvssHxaypXimglJJ0AFFELLWompOKgDjt0k5Rdg/TlkgRhZBBEopbzh2/Y5AvLNNFSZNVVXeedvUoam9Yw7egQNAMgBU9oVYAjzGGEAiLGGg8v3FMETJicFkcifo9O3tTY8vb9zd5CiCPuKII4744+BIQB9xxBFH/BHwsHDT8HrC9enpJclO1aIU34zMmnPXFXvFruvatt12Xd/HmDKOtWKcdYQkooBEZJzzZYLhZlcnc0KE2XQ2mc3CdAqAqkjNjNaaKPRqegZ+SqgUJa33/ux0tpjP66riLFU9ubi8sj6wQM5saOQZyShiYi7MpvDwlT/IZqHUMOcc2RA5771zLNK2rTUGEGOMMM52mHPm5L231hlDOfNms354eFCRPdn6D2lkHDVTex5jlPUIliJyRDiqfQn3kuiDPTzuCnDkbJ8ZU+CeEBwr2AHAaIg9VJobiuhoSXtGMgMrMVoDD6nJQ+l5xKH61jMGbDilkVccKMWh+twgEkMcT1VH1awwD3TjuHi0zXiqlR4MOAZLDxhqBemjNhxGwfVjy5T57jsm0cOx9ivqAZ8NAKBZlZXI1aEWq9vYtTG/6SIvLnRxfn5ydmEJ7gFAOMb+4fbLxGlxcj6dLiwQAu1gHdudxJ6sI+Ocr5rptK6rdrvabdfOGV81zWQ6q0/AgEouRcOs8YTYd7Hr+qqeTCfznKnr+8vTix9+dPrmbvnZqy93naix0nK5iYWGLrGDog8/lIcDqIg454wxXepUlQhKwjsAFpMN51zheUv3gwO1eiGgy00vfXVwdhEFACwOqqOnB45eNKqKSjrI6oeBYqDMyIeeoCWSMPbhQkY/SvQBEdFa66x7DDUcitXHDn9Axe655YNhMYQ9HhOr95bPjw4zOsZMyvkOeRcKKuez+sff/5P/5i//bOZ3lUOJfY5iyVvn0dkkkmJ0xnmD3XaV+y2ibLZt28r19SKEsNs8oMSz04VzdrVcffnFF+v17mSxOLm48k29vX17/3DHiWfz+enFhavc5v7+9ss3d7d3KjBfXJy9+Mg63K3ub1+9un/9qq6a+uLlMrANnz197BwK9/7J42uu8SvbYZTDiwNdOPfx5fmL08ks2AqpJl87mk3qpgmucs4Z520VgvfeWVsGCCFNJnVVVdaanIWZnR14XmsGdswYcs5474dOBWqscd555xCHgYaIIYQSHxIWInTegyqL5JSsM847ckZFOMfyUB5tavbpHohIoFgSQQgRrDMICMCiaK1xvjzujLUwGg4NUToiEeGUFYGs9ZMmtW3f9QjJEBljCY2KCKciEeYcAcQQWdLY95vt2gyeT1pMoqKxZfgjYoyxbdummdRVFaoq9X3OWVo3ZlooERnrhngwZ4IAmtpNGkLChGRscA5VOXa77aoMxFRksKKiknLq4q4IpaWaIJCwMrMIA4g1aIVju6uITGUBAXMfN9EQCXPf9+Pbbqh0l2JmLq5gzMw5ZxUBUGuoCNi3my0AhKoySMLctq333jsnwLHvu65jzgBI1jgXnA/OhWI+BlqCtboEJWtDHdBYAdMnCEl+/J3z1b/69LTC//M//Wqr0D/34viGnf9bHGrS0bc59v12uwvBz+fzk8UGi6dYSQVT4JxZREXKl4Yw74Pk5SMhxVjGJpbSHTbvGWrVvbgc0SMgKRYCukjhSzVsttYWK4xyXsOHwKFlkwKrsmpd+4vz+dxOELJKsZlSAOhS7lIGgOJ/Za0tH3CNd44IVXzwIYSqroxBJLTGOuecd9aSMWiMQUJDZMgCWjG+qib3bX8btz+5ytPuD31rjjjiiCOOKDgS0EccccQRfwRMTNv0Ws0mk+ksr1Pq80423HfctbnbceqFo0ru+76UQYspZxYXKrLWGLLWGOuQDKBD40PdGGuRMIRgjTUqdd34KqC1LKqC5CcMfr2LXRIuisQnQAD13p+dnp4sTuqqycxIJtQNIKGCMdYYpMIwGasAmlIpkcTMKgIjc1W8C5jZW0BEa4xzTkRA1ZiS4mtgtEJmzilHa60xxes2EpnCn+0dhL8p9IAgG3g6KXSzymDIAWAQeHAuQEAkIdrLf4bZ2ThDg2fs86BffTyrQw5aR/pYR24dqTibKOytKBAJCBAe7aRxPHMFGH0YcOAl3+Ge8dFjA4uweVyHSBUEgPZS12G/haxhLHwgjFwiFsdoPVCq73cMo9C7+FDDqK8e2edR/gp7erxc7l7wPZ7wqKEdmOw9xTmskzN3CcVOF1eXev9Z3Cy77XKz3hlAj+LraVXN5qfMHNuHvlutco4O0RtHxjfTOVqfkNr1CmRj0Thv29jPTxfWwHr1sF49YLv1zdRXNQBW1eT29rYKU2VIKS0WJ13bPcB6Nj85Pzt/9epV3q0+OZv+1fevPvvi5u1/vo9keCCV0Iw0kI7EBygUiXS54znnEIJzru97Vca9pJ6o8GIjhT3wyCKPQvjS3vt2GzpSySQYCejHhj5s4H0ffPwDcbTylJEoH4RniCAHoYkhZICoQ2+EUplqMCx4vKeHrhmPQtfDox90nmELHRX9QABCe3Z6tOEorj+KAgKffvLyX/yzP/n4cuZi6jfbftcRuNmsJqoALOfOkr+8nELcQlzXBhP4z9++urr+k6qeMnDMfTPzk2l4+/pXr9/cJMaTxfnLly9rX63vl69fv3l4uPvOp98/ubiwxkjcvf7lz16/vgnN/KNPv3f54XeJqN+u3vzy81/89Ccfvnh5fv0hzy9ze9uyHtQx+xZTUb9T4Dt68OEv5cFgEBzqaRVeLKYvT+dnEzdxUFtbW6wd1bWvah8q55x13tVVFUJw3jFLefrVTRW8I2OCApKZTBrnXOkyJZxJhqwla2wZIGiMc8Z5Vx52ososABpChQjMEmMPCtZaay0A9LEnIuuNDV5BOFlDpArMXMI/1rqSAaKiiGSISqE22Ov9URShOHWgCkgen2dawqXCyDkXuwzrvTcmpxj7VlgIyVhrrRXmPvbOWySMnIrZDwKkru+61hsLCjmnkqCTxjq0hWHvu444aR9y5/u+Z2bvvDEGEZm5SLDL5Yio9m0P2LatKpSkH+usdQ5Yck5d1yKAQRAR4SycVTRLTqlXVUTqrFdFVWBRAEEA6xBBYkzOOWtNHqoEKyHmnNu2HQO8WB78nEtJZB2i0UOEYLCSZ+Z21yqoc94Zo6ox9sX5CIBLIlTJ/yg5K85XznlUIRWDxCwx58xMxlSTCpBEISUlX89M+OGH89Repbb72c3m7aZPY2f9dRlVCk9W+LYOfB09tna73f393eXltXfOWgPw9DvGGECEwbccVawMtSLAWDtEzYuvGoCqlnEEIwGtYykCJASgkV2WooBWYRUiItbBCGrYdIhR4j6Gr6BZWRGcM9NpsKiFQC8fVDnloUMDpKwxs4qoSI5iCUHZddmHXPW5ZLVZa6y1zllnyFq0lowhY4yzHo1Hq+QnxjtRROBN+Lbe4iOOOOKIbzuOBPQRRxxxxB8BQZiNqbytvGsRus1m1e3a7brfbWK7BU6WtKpd+Z5GayogReOqyofKhYrIGOt9qIyrjKtt3ZCzUIo25QTtrhjyat8yS1aDJu7Wuy/f3nd9LHLfIYO+OPohAoD3/uTk5OTkpGmaxJw4J+bMGRANIpJRVckMmRUgM3POKcaUUrEXKJYC3nsAQERjLOe86/tiPbln4kqNJgUwxjhnKwylQUR0nHn+lqmRqjK6E9MBf1SmGaRCLKlQvcMiMoV1HmRi435G5e7hL2VXsF9yyMfo46xM98RiEbemkjxetqJCGqMSIT9Kj/euCIUxLKbDzAf158cTLmQPjQUVh2MXQwM84Atx4JULAz38YvDRahpUBbD4+kq5qvEKR/YZ9LEBRi+F/eYwEvWD8HnvCDF6ZeOYc/s4x3t0YCiXIxJzjgzNyQWZSMaQWQvz7ZvPOfYn5y+a0/PT6xd1Hbz3q+Ut57ReLZ2pZosz74MSzgG4j5xzH1vTYmaZz6bu9Kw4Qu52u7ubt4uTs7qZhIVLfd6u16mPzaQ++eDDt2++fHhYiuKLFy9PT08flg/Ybeekf/6di79/tfp8GTNj4aCNyTCyYGXSPbDPhb1iFhWRvu/64o4qos45M2QqKAAQptICZMqdFVUhouBDzpmZkYrjszjnRpJaxmKDOKrL9dFHdWz24daWwMYoR1bV4j1dnAFgn52gWmIO5TayAAOP3Rz3DuzDTp+ESPBAvAbwFdwMHYyJwk+UjoaPAwoG4RuogFycTP/se9/53ifXjpJzFHuo6jr4uq6rar64/fJGWSfzmZ9O2je/kNSnnHeJ59PTk8UidruuXYP2ly8ul7e3D6slGnN5dX390ceBaLNeLpdrIPvp9384nS8UcLNePbx9tdtuLq+vTy8/Or360DWT5f3dq59/try5OT09f/nhJ2Fxfp9wu9lst7vfOPr1TwlPomz7n96VhJcBrgiCAA5xbs3HlyefXJ6eTXzjNJBOKxcMGmQAzrnXNuVkOTsacz5KzERYoNWiuKyaejqdNtNmMpmEEHbbbd/H8kYwhqq6FuaUk/VOVfq+F1VjjA9BmXPOrK0hIqTMXPq8c85Yk3JWkJyzorLkGHvnHCGKSMpZRb2CiOacRcUaG0IYnDRy3ucdFG/iUrKPcy7jCIesBREZnHkks7N22k5TSjHGGKMqIJI1VlRS6qfThgy27a6EslwJ2eZMjQVQjrFEaoucmUWKuLh2TnPe9f36gVPOCDCpG2NIVVKMKgKIzjoiUy6qT6lrexYBGOynBRRFBtMdYVAxhCnGrt0N9vYICsgsfReLQ4P1RWStmXskqKsKistH2xKSd05Vc0593zNLqR+YMwsLoRlycAoHLeyss9YOeRyI1hgA6HhdSjUy5xgTM1d1UJWcMuAQ9k59TH1SAI69pt4Zyyx9TIqAxljvBotoMmg82jD11Y/+5Oz0pP4f/+f/b7V5qwA8JIq8J01nhL7b6b+tQCrpCOv1Cl+b+XzBkmPscmYWRWPKWmNoE6sqGGORqORJAaIpZTyIyjeAavFDN7r/NoDH5wEiAprx+2F4bXHOOcVChRflNQyfBHrwoQGEBkAi513fb7v2dDKpvHeutqMhmsjeV0yZuW07ALUGbfnc5MQsMeWYIhkkov19JFBjwDosjLT3gWwwVTNl27dJRIGM+Py3f/vf/+3f/oc/4L054ogjjjgC4EhAH3HEEUf84fEf/93f9jmKoc1Det2vdXvXtduYojUmeFeHUyhWDAbJWjTOWkPWG+tt8D4EHwI6j2SMMIoCJ9neCyiiCmeOXdpthBlUSGTX510iN7v+/Gc//fuf/KzdbAiBn55P+WwnY5q6zimt1+v1erPdtikLlyouiNYQqnLOgFRq2RSWSngkH8ukYPC7QEtWpFhQJiJyzqUUWbiUWzLGsOSSwBxCAIDY98vVcrVacebfcjK4F2zqwSSpcGeqoPy42qDs5bFqDsKTCeiB/BgP/vk46Xpk2qA4Iw8zOkVAGUWwox551IDSo2R6JLFL4x846YLuyb93Lw8G1fKBzHmkpscloxR2aAbdzxj3lBoORPA+1/ZQ5Tqejwx7emyWA4G5DozU47UNx9kT0I/M89B8A/9Z+EgAUEDh2PU5M7hQn5whinEu7bbr+/vd6s5aa73z/mwyOxUF46rN6i713fr+TjNXsxkFbz3OTk/a7bbbbdvNsplMU/BkXD2ZI5qcXnPfx912UlWzxel2s91u1sIJtaqb6eKU2y62bXf/8DCdTmmzanc7o+Z71/N/+enV5v/+/POHruPx/o2CrDKhHrl3lOKqMhZlEsllTp9ZStPsq/uN3QZhqByoCBBjHkRnCKAKAjmNac4wOGvsvV7KGnt2fwgwwOjGAo+9oSi1951zuBd6eIfH+IA+eokU1fR4jQBDB37aCZ/2yWeC2Ecp/Xj2o+B9YKZ1T2MiWAs//O6f/fjTj16eTUn6zXrdeGfJOR98MNv12xTXVTOv68Cxz7HbrldtTOia6+sXlbd3t2/7dtXUlGN3d3cnaE6vLi9efNQ09erm7Wr5oIgXLz6cTCYGtW8397dv375+U9eTxeWLxdUL20zbzerzn//9drWezs9evLhuXryMbb9d3q3evtk83KnKe2jY3xK/uz39foEHIYbDH5/9WTIoSoxQCcABeIDTKnxyeXJ9OjmtsMIYEGtHFtkSWkMIgkrB+aqqqqoKdWWsNWSss4YMADhrrCEgClWo6hqQ+pj6mHLOSFRVgZm5FBIAgMHcRngwzhcAICLrrAgXgw4avQByiioGlKmEUUWUxQKYwkkyO0QlhMwG0VpbXg6aEuc8PrZUVWOKAGCoGPrk7W6LAIhAgIN5v4gxxjvXS5LE3FthBuZipVRs/5lBAOKuFeauLxYAqFpqlPJ2uYGDWKaIFCdfa13hhlPKKcau65xz3vut20pOnCIRGiIiEtFBdCzCoiVIxixAoCqZc3CWCFNKCFqkrSnGvu+ssaXiIpFRwJwys6iC6cg665xZr5aiCieLnDnnVF4cqYslAldk4oTkCiMOuFdn74NZg3e2IhljrUEiBRUWGMJ7mZlVoaprBWDOAOC9r5tJqSYXYyKYGEQCENXMnJlHa26DAJyyKAiSWA3B2Fs2+QAAIABJREFUzhfnSfHyev5//KfP7re5TUCjs8O7o3H8IPh94BvKbH93Bx+e4EMFQSJDpIgY+z7lTM4Pr6FiHYOQcy6aAM65aAhijIYopgQKhKgiiGis2ceYdfRWKk98MmaMiQ6tK8ySuajdjbUYB/Z5fBTyKMYWVU0Ay7b/crkJjmLDTXBN8JVz1pgSWTVDzWad1Q5BEARKgFbdaFitOlQ6HPp/GT4pcxezaAJowTh0rVtzR6FPgLXLp5t6d+RAjjjiiCP+CDg+fI844ogj/tCIvg6x3SaXKK2WK699yjGL1tNZXTdVaHSva3UOrDPOGueN88ZgsVpkNKIiuccUNfW5a1UyKOfY5b5N3U6FUYVU121e94ir9OWrV7dfvo19X2qHFQ1tMbBUBFWwzi1mc06561fbza7dtVkGJaOqGEIsWcqAeqCRLERnEXOV5YUzs2RgnFsSGQDtY59zAkRjTRFqlZThumkQoe/79Xq9225/awX042RvJE0PKLPBzHjk7/brKSjuZT3jXp4KIHG0fj5YYfxhv+Y+zfeR1X30zNj/dyAoHZjD/dR31NmVln3Oge/PeE88wsEex9ndgd1BoSwPtcuPlPBeVvRIUB7g0bnhYMr4eJ7jEZ5oYx8tnp+07146PlDhBwcildh3fez6nBdNPcFTQ6Y3BDlxzu32AYkQtDk9byYniIbIbpa3uWvXfBPTLsxmJtSzk4WxLse4Wa8s4s4GGyrnw3R+2u5iv1v22/XW2qpuDFFT18I55xxjnMzmi7a9v7tbrVaz+axuJikxMLxc1H/zz16+unl42LabLrPiOxf/SFYc3rUiOgNEJAODshie4hlh++TvWNom7dttv9sSrXi8a487eySi94faV/rTMZ7x5G7s97InuR8X7HmvwvDhkzDCuM0zPlqf/TL2SX02fvb/lZ+9p4uTxV/+6Ls/+OR6Fkzctl3XLeYzRxYVU+zv3r6qqrquHaHsVsvtdvNw/4DWn55M5/PZbv2gcesgQ8ZXv/zlru0WZ1fn1y+rSdPttg/3d5zT7PTs7OUH/Waz3dyv7m/Wq5X19en1R7OzS/TVert9+/kv7m/eLE5OXnz40fnFBVZhd3OzfPtmc/dl7n7nCuhvBwf9GPx4+vP45/MeQIAWoEKdO/tyVn/nYnHS2CagQ6491t44g97ZEJyCOmfr0DR1UzWV96Ho+r0rlfeMM+SsIWOtd8ZaEem6LqdMxnjvjCHmzDknZjJkjJHEpZuVZ6UwEwIhsQhgSQXQEsTlFJWpsHIyFPdkhcF5Q5mRCAA5JyQsWmMVSSkXFxsAQEJV6bsOEK21hCbGuFuvjaFCzzHnzFlEgvfUNKnrQACZRcsRhyctkRHhGDsVFeYYU4lqMZeKDJBSRkTvfC4EcLGGByBKosrMMaYYU9/1dV0FnxGEU59j9M46a4wxqsAsOWctJV2NLeytQjHYYRRPBLHvEYAIQTTnzJkJCACZuRRxc9ZbIyKKCM4Y77y3QUQsOSUEgqqqACDnzMgASoR2TPvgnFQkhMpaW+x9yJBzXgtJL+Cdd94Vux8uZLkwc8byaWM9qzJnQ8aH0DQ1Z04xxdiXoq/CXB4wKWdhAVDrLAH0bceZWSVBxuDtdD5dzE5OJ5zav/vs/tVtm0FZYTQkfqfzP/74DSnjb44/BgcNRXuuiGiMtdapSE7JkClDj9Ngm75XDJRkHiQsZaVLNowhKkGCYjkFoAi0dxsDKG88InyiLi80cDGYKdzxnpsu9l/lfYeFMgbYdPFmtQvOxNhPvUlNyFXVhMohoiEEssZYSxg8gqhm1H1tCkQkRWAdumvxjRHRLJwT9ymlYuQBBKKxa6HyCoAqZ7f1xv3O7/URRxxxxBG/HkcC+ogjjjjiDw0E2kzP3HY5cZXFrrZWcCpoqnoSQu1cBYporKkqrAI4CyqICIS5b2PXbrp+vVr17c6oOFJLApxBsnLq+1ZyMqrOWYOYc1JVBNpud32XvKsBWhFQUGPQEDGLQBG2QF1VV1dXALhZ72JMfR+TSPEHYGYCJUIik5iFdbCAGE0FCYmHTNiRlpZiHIwxRiKMMZaKRswse7mvqohsNpvig9G2bdqnPD+KjP8hE7NiylHqpRcCBYnocK6nj0zx+O/n+xj4WxzJGd3zfM83UzhcayRxR+ZVR+YPx9N55JL3F3tQ+e2QND743+NhaSg890juKaCOklcYawo+3RrGhXhgLfJswV6tOnpCv9MoT3nr/U16Tkg+MrjPOHCLEPt2t16tHx4uq1moJihIiE0VNvf3q9W671+rChobmmlVT8iQ925z92XfrtfL+67vzy6vQ7Ows5kRcaCb1Qpw7RNDA7aZnp5f3HO/Xj503etd24W6aZpJSnG3293e3FxdX08mTd91Xd91XdfUDQLFmADNjz4+/fz71zfrdrm7X0fRd1t9FPgeQPftvW+Jg8jEu7Pc5zq8p/7Kj/3lsFGHG/nIJr+HEn7eDQ+DJjju8evG06FP96Hu9d2reDJIH4/ydUuHs64n0x997zs//u7HL06nmNbb5bKuG+u8QUxdu1pu2r47vbwMlUtxt90sb25u+ra9enl+cXERY7+6exMMGGvX2/UXX7y6fPnR+fV13TTb5XL18JCYFyeLk8sLDD49xNdvXi/vb+tQffr9H80ursiE5WrzxRe/+uKzn5+fn3/48cen5xcAkNer1d2X64cbjm1w/2V+GL9XGzrgSaRrCHepRQoIFeIH57OPzmZzDzNP08rV3lSegiNnjQ++ripAMMY4G0II3lXe+VIB1RbfXyRnnXPOlnKdOXMuMkYxCJqx2+76rospqqp11jtXyCYkqqraOcucc04pRgAARAFJKYGCNQZVi815n/q+73KOgGrMYC9giESBVUV0kBsbg0SIlHMuVjbGWkKIMe7rDTJzTKmuKkXabtZd18WUiMBau3Qup6wChMYYg2RENcaUUnLOsXDfx2nTOOtyzjHFnLO1xjnvnOOcVJVIU5K+TzHG2Ww6mUx3u23OWQVV0BoX5jUAMAtzMgDeexDJmVVlPj+xxu3alkWByBiTmVNi40wIvm5qYRbJwlw8cor8HFS98wDQ91EErHWLxUJVUuqLgJmIXn7wcXEHUlEkrKqKmWMfAUqducEHn4hyTszZe2+IECCmhIihqlJKMaYUc5FvxxQzM4sUGxYWaZrGh9D1sVRcnk4mzjsEMBZCVVtjVJQ5xz4qQKkkMT5uRYWLxbYoZ03gnKtsM6nrupk2zb//n/6v9fKnuwxxiBN+DSWMX7fw24EykDEzxxhF1TrbTJrNdkPMxhgqJSOQy8fQIHwnIhpCAQCAiCrDu7t86Y2hbBBhPXjNDXJjlGengKqRI2YggsHZadidoiIOhT4BAAxAn3i57Txpu5YG+SHYaV1N66bxvgq+8q4K1jtrvSUDhOCdM4QKoDI8kZx1xhTLZ2uItCQdWFvqkbCIIikSo0vU/PL2oUNzx67m31rrcMQRRxxxxG+P/zK/s4844ogj/phAcpMkJtSL+cJEVzkUBEHyobIuGBsAQIU19Zx3CgIqLDnllPouxj7GmPosKYkwExhSkKGAmCoR1eQ8jbKoAG7C7m5LaN7e3W9izONZPDIOCOCsqaswnU5Tyjnn6WRKzrOWAn4AACAMoIDIo7JmPw8prJWIAKAhGvwKRAjJGDNqnMR7X9wYABGJigFu8Y8u2bg73Ok35Zu/wVqPbJg8srwqyk+olgNODh//+r4DHvB5j4Lfg8ONFscHO9JHeesgFd7PDw+YStwz4Lrf6IkF9fCfDg4Wj7Lr/TkcENAAY4L84boH8mMdhbB6SGLi/vCIOhDQo5D6/e3yhIB+9sPzlcYG3nOrDJD6vl0t71798ipc2pPT0MycCxK3KSus13G3TruqfbixBH46qyZTtMCQ+rc977bY7lZv3zpbV5PZfL5ABRFdP9xx3DmDNJ2eXZx5oyp8d3e3Xj/4uqrqBsD0/fL+7qYJwYeqaurNbvvZL37xySefNFWFAm3sF/P6v/ru9Zvl9m7d/ucv1vmJfhie8HRPKGl458eDy36+TJ9Rus8jGU8b+z27fPzXM6X1V4dtnhHj79vqyYV83RB7tuiQn4Sn/eC57ttbe31x8t/+13/16QfX2m6363tP9vT0SkXW2/vd8q6LaXr+MiyuBHi3u12vbtvt7vry+vLyWkRuXn8RNBnR7bZd7frv/+DHpy+uvfXdZrV8e3tzd/fixQezi2vrXX/zxfLtq8+/+ByNv3z5cn7+AVrLOd7dvH71q18sLk4//d73ppcvQLT/8vX9l798/dlPWWl+tjg5OyV6PQ6i3xS/OxnjPwo878Djk00J1IDUzl3U4WI+O5tPT6ahsugIg7EWARgEVZIkYgDoOKa4csGHunLOgoKIkBn4L+esddZZqyAijDRUhR2s9GmQMBtTivnZ8ophkbqunLWqknNmziXpYyzjiQZL3BYQse12Xdcag4XzHgsSmMySVQGQhYXVeWeNRaKxuK4Wzg4RhIeUnfIGQyBCSllFCMAAAAtqLBFdyCqeLAFmUTDWGUuGlMUIuqquQoWIfd/nnIL3xTU++BoAg/MxxcJZV1UVvAcBEUFCYQFEa1x5ORCys2gItutVMVKYzRfWeV/XCojGOu9YtHDTxplQVeXtZAiZszBb54gQVJ2zoBgTiyiRqetGJMfYA4KhobAbIrFwcZBGQhI1gVmyqtZEpd0ANeXEOReLbRW1JiqAWleqEatLxli0BpBQxIBaa1VBUwQf1HoCcsaaup5MpwjYtm35kLFkUs4S0ZHREvgmRAARzZyUwZAnUFBFTsXmi1Auald/+uFm2Uum//3vPr/dtO/WFx3Dwv+UgDBEBlLs4zSE8/PzdteKqnW+BBKcteXtQXvD5aFvD6YzVBHCkGEAw4sBtVSnGN86h7Uhnh4eQZW5lLvWA8+yQzwaSouqIvl6Eqw4TUQqDH2fJGsf09aQt8Y6Q4YAFVArH5yzdv84MEYABNSAWgRjhjM3CNaSWijDE5DIea0mvfRv1nGSKsb4e7wJRxxxxBFHfAWOBPQRRxxxxB8aBpRAp/P5dH5iufYWGSSrGGuJLJJXVO22cX2f+zXnDgFi7Npul5hZWEStCw5NZi72vwqgapSs9bULlQ+1cdY5XzeNCxMGH79YZvh/394sexnoIi3TawAARcTgXV2Hqqrb9iGnNJ1MqslUiHJmMsY5wzmpsCrIyDcOU/2xylBRQhuiIjpRUUNkrSGilNJ2u3POFZNN65yxtkyyy8yZmbuu26zWv0krPp0zfr106UCXqnpA4T7Z1bvbP6fPvnKTZ0n2o40FACjQ+3ajB3soXrxFIox7v4zHAzyy0o97PuBBD+XSxeii0MHvCnX3uyh7kL1AeTilsTcMBDQ+MyP5iuz8/fzznaPhOzepMNylEl7OOcUectzev60MTWZnzgd0lHM6iX23XoLy3c2bXdcurl7Mzs6reqKaOce1aNzstnnd559PF2fNbB6a+vTiglB22816/YAuAIj1bnZymkRiStvt1rm1IdvUDed+vV6fh2o6mbZd18d+vXxoQpNT3q6Xm+3ycrL4l396eXe/vntY3eyY39OKj6Kw8aZ8E3wlAf3N8N71n3D/xZ5liHocHvDrCZbH3vbV4ZdnquzHv+DTa9GnQ/FJ/0GA09PZn/3g07/88Q9qq91qbVQvzi6nk3nXbREwVGG6WEzOLlGw3W7X9w+b5eri4vrs8qWzrt9uMMfdbqMawbiT04vzi0sQfri7WS037S56V03PLxBxe3vTrm7evvmimUzOrz988dHH4H27Wn3++S9u725ns9mHH35cn5xIt9ve3t6/+vz+7Rd1XU8mi5XNzfTufQ7s/wTwXg378/v6Tk85vNEAoICKCgbAIcyCvzpZLJpmEkIdPEnSnMVQzArKZCja5LosqrHv15uV8zZUoZhscM5UjIcRjSFryZqhfpox5Jy11pasGmvJe+9DCN6XkrYAmlKOMXrvrTWIqCrFxDxnZmZrLSGiavHHV4Wub1Pq67q2jhA1pSwigJRYsioSARKh8cFbY3Fw9lccie/gg6rEnDkxIjnnUxZEQBNc5Z3qoQmBKghgCMEY28VkrPXeK2jOHFKq6rqqKu986LucY3CBEEE0VIAABsml5H0uRgeZBcl5R855AC3CTmOMsyZ4W9XWWLi/vem7npCqSWOtq0WRLFnrQ6UAiXPsW1Ex1hrjjLHOWc5ZMvvgkUCViQiAWECVCrWbc1TvQdVaF6pQRoQZ7K45poQE5EKKPRGGuipGzKKCZNFmJWIFAVFPItKrGuvJobUeABkRYCh2Z6wV1dRSQhJRNNY5b60NVc3M2kfy3jiLgKqixljvAaC4FQOAMgOIgqAbqtBpsgqASJBiZdzJyelf/+hTovD2btPFzDGNodfh1apAT4OK33Yuenxxqyrnvmtn89np6en93V0fe2OH5APvnl+mWKuqVKpflhEECKpECAAigjiUki6BobLVWB3hGQENUIr0qgCIclZhKN+bxYBj2HhoblFEstPZYu6x0ugkG1UEyAK5Z9BoCIlIUVlFlL1z3rmSXVENjwUmQmsoeGZ2BEAExqCxaAyawU6MKusx4MvT+UN721OH+jV1KY844ogjjvh94UhAH3HEEUf8QfEf/93fgma2zlmHaKwPAKKSRDm3SVgkq3KS2HK7lNyqJELInBXAWUNCKTMzA4IxdjqbTGdTE2q0XslRNUHniSyKADMIY1UlcT/5xS9//vkXSQAACIEBRVWUi7KMCEMIVaidczHG9XqzWi7VOnIuZi6pyin2quKcyaKiSsWqeFTq4pioWeYn1lrUseqaKABYa4uUDGCosEREIYRQVUQY+9h13e9n5vd8SvmcHvsKHeqjivng13c478MfhnJu7/C0h1Lpdy/xkD882BTHPT5lhhQB94X8Di5tL8h+lEI/Ubw+YwkPjvHuD0/Nmp+c836Fr7qa57+WvnE4vS/zTy2/IwJp6lbbtYh0qZmf1LNZNTkBRR/8brXc3S+72AsAEi3OzpyrZicXhG5L9+1us9ut0SAZbKbz6ck8c0qqfYyb9T0SV6EywTezBa+WKcbtdl1Xdd1UzeTlzc3terOpJ81sOs2xT30fARGAQHa77SL4Pz2v/+LTq1/drDY/u9ml0oW/ut2+ui2+Anrw5zfEO2T+86XweGMORdtPNnraB97t+Y/Lnxuhv3N0fHoV7zLU70HTVN/704//5i9//J3rE16/VeVqUoemTn3Xbjd9F52vTs4uXFXFrt/cP+xW20k1vXj58WQyhdzzbtNvV9vdtqqr+cn59PSSANvdZrNe9pH9ZHaxOG2Cj9vl+vbL1fI29fny5YdXVy+bqpJ+e/vm8/ubG+fDyw8/Pju/ssYtv/z87otfbpb3gjCdn7jFRcitotGvZuK/zTiMmT32lMLB8Hu3GNYp8SiB4TlT3BvobDK5mE0Xkxpy2ix73SFpJmBnAEFB1VrjvA8hlEcKEiXOaZfJGGtscX8u9BaraBZmcM5Ya0SHzBhjTHnK5ZxVVZgLAb1PvikhTEQ0pjg429Izi0GHNYYIVTWlHKo6VJUPjghUxQcCQFFQg4AoCrbYgFiHgMxinSFCBMiZAbRuagRk5hgjIHkXyruU0BIZMtZYYwwhGVUFIDTG+YBIm12XmRWhODLHPqaUNwk82j7Zrku8aUEKXSh93+92276PnBkAYowxJWdtXTdN0xSj5KqqhIUQZ7Pm5GQ6X0z9yYsKEVSFGYnqqi7O8caYzBm1I+cNgvOuVCns+mSt8U1wzopySsqiIiyKREho0FprDFrPnIgIjc05iwgSWR8sIqVYxLLeEBHawdMZEMlVzgP0sWdmMMZXlYh0bauAxthgXSHWg62MtT74lHJM0XlfVKulQrG1tthq+7oiQ4ogqsZYCGQM4VjWVEQwExCQULnpgKqYVZQAWbqYYo65MdV3P7z47/7VD5y3/9vf/RIAeIhE778F9oPi1z/E/pGjFEAehczQtm3f96GuMnMfkxGgfS1c2FfUxbFOJgFAqRFtnSsEtDFUnDdKpUHmXKzSCx89dJxnLwsdyhAoDMWfFYBTBBF453NCFWKWNkrMCsE6VzWGvEFb6h8qGILynBCArMVvPYtI18e+68ozyVpy1gZn67qq69pb47wN3njvwBk0xYRN+r7zIVfOWSVRIaV/86//9f/wb//tH+bWHHHEEUccUXAkoI844ogj/qDIYG2/NXZeOwPcdX2XYyeQFTjHKDFLyiAsOabUKTCiGmMz2IzoQ1U5N7FOkIDIWNdMmrrojxAVsGPmbpsVjCoyx3bH6806mV998cXN/UNSUMInGadYGE2sm0moqpw5pbRrd/f39+iDr+vMZaapCAoqux0DEtBQdmbgCMZS6SVD0xhDiCJa5jZDujQzgDKPrh6jgqaw1THGko+sJYG5LBrP8RtNBwtX/OuUiwd2GL9m59/goDqSzmXm+n4V8K/f0zu08J77frrLQ5Hqe7W0g14Pnq+Awwn+GqXuvl/sSw++d/Wvv5x3Wcsn5gyHvKax1oegzLnd7lKSPklONgTjqnqOQNClpKtV5rR6uBUVg+Ank2aycK62JuQvX+U2M/dduwKEZvKini2yoizvd9s1oORmWtWTZjpLibebddtuQdnNT05OzzfbdrXZJObpdLKYL+5vb/p+552bT2uCrHF3GqY/+vjsF29ffPZ283rZ9lmeXtQ/CL/J9l8TP9jjufz+Ocv8253vr9/wN9s1Inzw4uov/vkP/+LH33Wy2+0eppO6nk2zcurabrcREWNr6yrNcftwt7l/QKar65ezk3NS6dtV3C23q3sIVXN2Nbu49iG0N2/Xm1VOuZpMZ2dX88WJbu7bh9vt6iH2ab44u7p8MZtMUrdbvn1zd/ulD/7i6oPr6w+M9+1q+XDzZvXwpQgvLq7rxbnWC3mbNm3/D/Od/8eOfRlNfDo4n4fbnmD/TFYCdYgTa8+aeh68FRaOkZmyOqOWSm1AJQJDBgwoqbXWOReCBxoOaa3z3hljiwEAgFJ5qyAgKiE6a5z3OJZ0ddYaaxGwZNuoirXWew+IUkhhADBUwpk6kKFoy2tR1aZkDFprjEERzpyKPZRxHql40gIZY40ZCXmwroRLIaekAJPJBEBjSj5FRPKhKo5TzlVoPJI1ZIFQATbbdrNtt7uNwC4mvl+u1tvtruuNcywa+7jd9pzZ+/LWi12ftVREFIkx7nZtzlmYETGmlDM750IIxXYZEb33khkRmro6P5tdnM/ns8l0UjchWMI6+JNFqLx31qgSgyrZUJW3NPR9L8JkjLXG+aIxRxbJiQHROQcAAASIiMYSGUsAIMWPBrE4HhARIOacWcQZg4iAyplV1ZWlAEQECIRkrEXm0eYBBg/iEl2w1hrDOVtEUwUQKVUlCRFFRTIUgrukBYkiqjNEhUxUGD1ShLD4XRvmnHJEVSJyxig7jUk4O+KrRfibP/8U0GSGn7+6edi2GUCHoEoJQz9G7b763fctAGIpeiGgKiLr9Xoym80WcwBQlZxT+Q5gFhg9oItQgIgQQJgBAJByzqVIxF5GUDQGwlwco/dfPirPjdNUtZRTBlARFhbVg8+ux3XLJ4dm0ZilT5zYgTWlf3prUJRADYEhJAJFELUsSdQNmXfCJQ0PQQGYRfteRXJnjCE0hhBLVIOIDBlDxvktQJhtYkyIZzxbw2+UdXfEEUccccTvAEcC+ogjjjjiD4qsmLGagEyC2W1X6+XdZn1vDThHHKOmBFkMEat2Oaux5Jw1dUbIoL45qU9OT0/PwFm0RkuFcc7QbjV1ktrVmze7zRokV8ETwnaz7RLd7eDm1avNdpcAoFC/wkUpAygqCECTyTRUddf1Kaa+6+/u70yo6pwVKeecUppOGhVerZchVM4HgEHj4pwvfn/ll5xzYcNTTIbIOTdmaKq1FgCZWYuSF1FFmLmu65TSer2OfaeS9xTAN6GJn67yjkfEV614gKdax0f69teTb0/F1E8Wjjzrfsr1OEEbNvwa8u6pscUwG9Zni0fongcsvBLunRVHPnlQqD+u+rya3QH1PP6rcEKjGcgz6EhlP3MqeFciWy7gfdJZBQDn3GQyJbIgiMqc2t363jbN5OTUWGOqxjWzerZT5t129+XrL2Lff+d7P2gWJ6Z2nIWWD0564bjdrLouTZpZM1uQcSml9cPD6mGJaOt61jRTZyvOsny4SX1n0NT17IOPPv7pT396d3dvrWnqxlq3Xq1B3IsXV80k3N7cGMxX8+pHH5//P7+43fX5btvJN+la3xS/VmD7VdT/+znosce8K2QGgAP/870+/iBicrjBwZrPBsn7PSmesQ4HKz7XEiJg8O7HP/zuX/+LH358Mbt78zPIsbk89SF0u41Rtc5Vrg511XdRuu7NF7/Kkc9Pr04vrhQ0pt16fXf/cBtT/8mn31+8+MAQdsvbh+X9ertt5idnF1eTk9Pd8qF7uHt4eIiJF6eX55fX1WzGwrd3Nz/76U/ns/kHH35ycnFFzuS4e/XZT7bLG0E2lT9/8UGYnqw73m02y/s70WcG0F8/VL9NwIMMeBo83n9NRsMIRVACsAATohNnT+u6Jsq7HVoQp2KArA3eGAPWorXUTGofvHG2ruu6qquq8lUw1jAzIllrisdz8d8outeu7/q+q6vKWFsyb4rLazOZhBBSSrvdrt1tAbSqq9lshkgxxoeHhz5GBKgW87puvPcpJZH9TVQR8d5570Alxb7rWxEJ3i9OToogt9CmzJJzRiTvHBnch1QRcTqdZs7QbY03ZGxV1yII5Kp6quBErAIl5j7GL1cPv/j89c/+/ufbtl9udq/f3rx5e3v3sEbnRCDGvNsmZvUemTUlbTOIPI6Wb/6YQYDzRXV9MTk7mV+dn728vrg4mV+dLq4v8vlitpg23pIBQcDppDEGUmpFskhuGu89WYuGAJVSBKulAAAgAElEQVSYLKMask0zTTnlnEt5OER0zotwSglUjTEhhPLWLhSkiDjnEDTFmGNS0OAciIiyIXBkjTEiIirGEAGgaillDGRUFIS5F43JAFRVkMzFmFuZmRMAE2Hx/S2ZVVQoRQUtTkx9X0TZKmLIVNa1KcddBwg+uBAqwBqMTVFAZGrgn3//O5PJvK7rf/8f/tdu13WgjPuyCu/09W98F/6xocSgyw1kkeVy2UynV9fXZaClzKKirCllQDTGcPkeVC020Nx1QASDkB/2eWwH+x+e8yqMhMZafUcAXVBCBcIinFUyjpbR5fNOD143opBY28h95mQxZXFEoEiGDAABG1RCGKlyY0NVdo5UHiEU+y723egP00mvOXPsc9d3MWUAct47H9B6N91hPWspJGte0aupnf2ebsQRRxxxxBFfhSMBfcQRRxzxB0UUFEDbtjc3X4JE4ajCSVgYQZgAjbFkjbE2eB+mMzeZkQvCoElsPbHWpswcU8qp71tOEThbZZDEuX3z5lXq20lVpX4HqqiakmlbWa2327YvyZCKaNAW/z1EAlREnE5ni8XJZDZVIlatm4ZcKMcCAGMM56zKhmhgsEUKS9X3PTPnnGh0wWRhQhomkpyZBRGMscP0UjWLiKo1JnNOMaWchCWlJApI9Jz8+R3iHzitxP3/cU8P6+H0bJQOv5+4fXIiz+a9ewuF0V/jKzWYj8x2oQz35NFYC2hPMeozXlLhgH7ec9LvVUYfFB7cF1WEx70cXsWestfHy34m4f4KOO9mp6cv/vQ6ffkTjS0Lc7t+++oz0TQ7u6gmE+v94vRku3x4+/pVd3Nz8/YVGfrg4z+dLs58mJxffZDj5ObNq269Ncrbh2UItQGcTxb+pXm4u20f1kbQXtBkdnp5fd13m91qtVktq2Y+AVzMF4ZovdzmrKfnl4jcblf3y+VkNuszb+4fXDX/wcdXf/391cNm08V+G38HstixWd9t098w2gJP4hR7lvdRJf8Y8MCv4K3fo1V/fmDc66/f3eadzYebPh7t6cggQ3/yyYd/9eff/+7LkyA7DK4+mViE3Peg2KWUEjtXeeNR8vLhNnVd1ZxOzq+0bmL7/7P3ns2SJFeW2BXuHhGpnyzZYjAzaOwIzM7u2tKMth/40/Cv+IUfSCONpHG5Rs4uMQKiG93VpZ5KHcLFvfzgkfnylQAas4OeATZPV9d7FRmREeHuIfzcc8+9/fbVl1cvv4EYf/DHX0zPnjBwvZrPb6/rpi4Gs9mjT4eziXbr6NdX11fRp+HotBrPyvFJ225vbm826/r55z8ajyfj0xNb2G41f/Gzn3779VeuKk8uLmdnl6YYEdB28XZ1/S3EBjU7lb6Xm/Duif/+8VS5Oh8CIKpFZEKfktzfsA7O6GEehIISACMO2ZwNB2ejoQMwoEVpS0eFA2dhUNrSGcNQlm5QFa5yrrDWOSRiY4xzRVWWZQmIhERMTFkRS9YZwyyqAxmoqnUWAGJK1hjrXOEcIKaUgqRyOJicTFWViaxzkoSdKwbDTLkR57qDSNYiACGpiuZaapRJs+iYes9iJEAgJmJAwqyxBcSc1oOUA3EKQIrYBAFmHoxR1VhXDMbbut1suld3t2+u5m/e3s0Xq/liNV+ububNfFkv19uQUoip7tq2822IESQpiEiMCqqcQBWSYMwlAHYXm0Ku6fCbQQA3TdhebV7Nu+rVcvjzV5Wzw8JNK3c6cbNRMayKy/OTJ4/OT6aD0bCsKkcI1rhOTWgTiM9uJarYta2INnUNAFljTkjGclkUqtr5LvuchK4jQlDIj3IkghSZyRBSYVVVY0gpxRSSiILuOUdQSNn+A/pbBSLFGLuujTEhYuFcijHGqKIpJZEE2nuwWGuYGEC97zrvU+p9w7IddUzZIowJOaUUYlCNxnBRlYqsSKpIQADdtm440p88O/+3f/45Mv70qzdJ7x9u78Zkf2+hB/UnACC3mLXWWstsYkr5sU3GMLExnPp60bsxR5yboa/8+fG9EDMASPpo3WgRAe3V0KAASofxcoD720tSaGOaL9dF8lhyTVJZUxWusqYwaBBKZ4rSMDMgZbMXzQFhFRRBxFw5M78V7dy9UQXzzpOqqEYR7wWLCqrKe4yKg8m0adv/2hY/4ogjjjjit8SRgD7iiCOO+F4RJRHGtvEbAwxBxCsoIRMZtmzYOmvJGHLGFtaUJbtSkSGKoqim1IXofdPUTVN3bS0pgiRnGDTF2AXvVVQBfUwIUFWDqigLSZvGr+om9dzUPcnZzwkIq8GgLCsAElFmPjk9VWJkE1LvwYEqqslay8YiUZ6CAoJItuYkwl2eLQAAcLYIlJRSAkBj8uNGRYREBJSZWZiZmbiLnfdekhzOT/bTmt+GkHsHH9z0ASX3QdX0Bxbhw98OD+4hdfMdSSm9p4AfbPi+h/THtn6oYu233lGGenho/XLdz/gOz+eD08ePnMx7q+6KCh2y3N9pGo+ExnJRldPTc3axW1w3m5X3Xdwubt+qgEzPHxXVwBXWh1CNxz50zWa7Wtxa60RgMDkpq0EyUA3rrvb1trG8jklGk9loMBy6MnZhGe/q9RqRgO1kNDk9uSClEOLV1dW54mAwANX53V2zrQdFURRV1zabTa1IxhZJoooMC/m3P3z8Zr5cbH19U/+TREZ2XfAxDvqfmtNUhYemOx/a+8Ex3I+OB0P8u/brh8DMk9Hgv/vrv/iLHzw7LTE2awAYj6dlWXSd36y2q9X6ydOn4+EAJGxX9fxuMZ3Npo+eFaPh7c3b67e/WC9uykF1fnI5O73UBKvNajG/3azX5XBw9uRZVQ267Xq9eHPz9u2m9ufnjy8vnxhDCLBcLm9ubkXp2WcXg+HIOl4vbt6++OVq8VY1jGePL548G89ODZjrt29u374KzbZ0Bt+5Mv/QoADIgIbQIoaDqNm7ndynyO8/U0c8LYqTweCkGjhNBUPlTFlQUWDhYFgVVWGNoeGgHAwrY40tjHUuqRKxc4W1NhsvZAltLgyARNYyE6kqkiNGQFRVq5rr1ho2KcUkSkxFVQwHw5xwQ0TCwmqQkJBoZ/ckoqJCiIY4lzFk5uzjkONpROisRcD9U2zf2UQMPXvVx24USRAjkKIB5m3Ttps2XLfXN4vrm8XV9fLVq+uXr69u54v5YrlYrde1tl7T/jrH3uohah+zzZcSJtg1em5zPLzefv3wy6FFVAgh1T4hdASQ/1iEgmA8oFFlBqV7dHn+/Onj8bCcjgens8FkVE1G1WRYFYYsgSEwREwUOq8pZjcUVc0xYyJsnct+GCkmUW0py5E1pUTE1hoApf7dhXtfjhRT9uhVUZV9wCOllGJMKdt5ATN7H7bbDSggkWUTU0wxgmYGXLAnoKmvM0nQNE1d1znUbYzJEW7vQ44lpJhy+UTQmMvaCRkgy9aVxjBxF5JQObKDH3563nTtzWJ5s+k2PvWm5geN/90Sqf6lQnOh6D70mFISEWauympQVTFFQCQCRLLGGDY+hOy3LlnZvivpQYSqoOndh96O4EY2BNnK4yPh8vwqqD0Dnc098J0XvPwnAYQkddvVBodoRENk9G3nnSmYGKEsbOmtKxgIFNXEZEx2XUckRIV8m2BEZuS8mBiRiRgBk6YQgw/R+4huQMNxXHmNYVu3lTnSIEccccQR3zeOd94jjjjiiO8ViBJTAkkS1YcuSceGXDkeDqZFOXDVwA2GaBlIITXNZlXf3ogPEoKEGLqOAMvS3d3dbustMTITMwVjsnRoNj0hNqIQQiQ2k7PzYnxmt1L/j/9psakjAGs/RclKq5w9iYjOWgBcrzfBx6Konp2eB5EgQmwAULJwS4UIFCAmybabu3I0uE/MhCyhSgkUsk1gpgAAwFqLCN4HwF4cZZittW3bXl9fv337JsUIB04Hv/Us8P1s2neYNwRVVEC6Z3v3s/3vRq/pO8zcQzJ6t8v71T+yPH+oh+f6258tPCCPH+ie9hTG7n98bxc78dc7TPW7x/7+Cb67ynuHrh86kHeBCKIaYwIyk9ML7xiY/N2N+LZZ3WXP0MnpObmCXFFNpgrKRO1ms7y7UtFZiuVwjGQn03MQWt/Nm7brQmCi0trClaPxOCW/Xi83q5UtqmFZDUczUa7r7XazbrZrZ7lwbjio1uvV/DaWVTmenm3rzXpTT8YTZ7Vpu9RtP7+c/Plnly9utjebsGzjRxrit0Tf7h9h9/XBeu9teDB238Fez/fuF7/PD3xktH/MjAEPx9KHjnnvobpn1HpWDRFxUJWfP3/yb/78Tz67HDtpm3pbDieuGjNpDOu2qZ0rhtMZsyxv766u3gjAZDYbDYvWr26uvtmsFsPhYDY5nY7PmMumbRe3d6v1lt3g9OLZaDz2XbO4eX17/XKxXA7HF8PJrBwMJLSL25u727skMJlOi6qyg7Jd31y/+urq1dcW9fzy8eWjZ5PpqWXTrBbz65dts7FFMRyNv4vjyO8vFLLPMjEA9zfN/cV+n+XRr3ufYgEGcWD4dDSeFmVFWBpbGiisWqvOaOl4WPJw4JyzZVVWZQmEuZ4ZAzKbsixB1betWJvjjvlrmaGLgQhd4RgJVduuZeaiKJlQUqzbBhGJaTgoDZsUQ/AeEY2xxrCI1vUWEQ2boiitYRFt25BAjYUUvMSkhokQCRghxtS2XbLWGsNsVDUlTSmp3IfvRPKVjoiQkIQtmDKiabx89e3yF19+87Off/Wrb169en03n3ddSD3tqppUWoGkwAfNLQoCQLi/DWM6IL0REB+aOX0XAfT+9iG7v3OtyKBQJ1hvxNQBMfzdm5Z++hoRRyWej+nJxcmj85PL2fjJ+ezx6XRU2cpyYZAlMYghTTFJSogUg/ehkyTW2eFwCAAikks+Zk+SbI0Sgk8xxBTLqrLWalJkQqaoKgqikJKk7GwSY4wxpf49wRgTY6jrJo8EIsx1Dp0pMlmpqoTIBo3piAlRu67tug4ArLHMFhREUAVyeYrORyK0lhiha/1qvVk3ISJVg9F4WFaFTUm7CF74YnL+Z5+fr1d3/+WrW3+zjf0TSwHo/Zvy7xu0Dwpnex3Mra1IOJlOfAit70SUiJnYWGOMcT6ISC7jkXL0RjX7p6tILoaZsX+7AwAiJOIcith5rL2LPQEtMcXgfdu+78Yl0HuGCKAqsbFFWXIATbFrffR+C4CamIgNsiUyRIZdUVRVNRoPq8o5NgCqyAAEBEjIxEzAmNn0BCAEyRgpGXhYmGpgxxOxrZ+vBuha/Sd6ph9xxBFHHPGdcSSgjzjiiCO+VzhDYmnmRhcnI8GpsBKRRWvJEVoFaurGRx9TB9L6ZhOarYZACgwo3itCgGAIqsIpqDFsLRs2xjrrCmsLLAp1ZQJEpIKY3BC6rvGh9QF2jKD0LKGKAAIyoqTou7be2m29retayNS+64IvyoECxBhAFUCJgNlm/+jUW2zEnnxCJERmjjGmmHL9l72kBgBijFkTnWvf5HL2KaUQwjvlB3+HeMjE/qb9HdprvL9Q312Chz8OCNzvQmc92PbXYs/1PzD93f16LzA6VHHqjiJ8Zzfap6x+gCj+r89Hfu8MEe4LHAJ0nV+sVqvN5uR8MDw5F0QfAkiMXduu5gsASbGYnJqiGE5PDDOqQorNZnt388oHf3b5tBiOB+OZdQOm4u7tG42hWS8toY6m1aBSnIUUtpttu92sVys1RTU5YVehim+b9QrGo8lsOvXtdn53c/74yez0FI1dfbuyJ64sGFS323pg4QdPT7643rxcNJtXC/knUcf1IYEHbfOxNvswDa3vrLPb8oMH9460+n4IfHgIvnskeFA78nA4H5qz7DO4D0toAoCqMeZsNv3xv/rjH33+aOw0tbWKDMcnim5bL7brJWg8v3xiC9tu53fzq7vl7bPHz11Z+Ga1Wt5sVm+t4fPzy9HwBNWGkLar1Xa9RrKz88dnjz+JvlnNb26u36yXS2vd9PTUlYXvmmZ19/rlqy7K7OT84vETNty227u3387fvuia9ejiyZNPfjCZXRDSZrm4e/lVaFZlVY1OXDlaHjjb/GECAS0RoSaQg9vFh1ZUANBsRzIqilk1GDpbWZOJy9JhWVBZQllgYaksnDWGCA2ztQ6y8YViUZauKKwxmauyzmXrDeeKXNQOUYmQGDNhVZVF5jfbthUVaywx5TCnSkIEa5gou0gjApaFQ8Ceb1JkhEFpQRRUCkNKoABEgISiyRBy4RCBUJlUkookkCQCooDIigRAriiB2Ic4X22vlotvb3/26nrx+nrx9npzfbO8vp0vVuvVtm3ahEiIFPtEIVBkRYiS9s2qB4HQ3Z06V4oD2AV9PhJregcfiP+8c13mzZKqT4qImpL6CADbDtYN3G3kmzfbYemmg/JkWJ6N6cn55JMn54/PT8dVEZOnvfdCDi0D5PByjL7ruu12WxRFURQiqin6FImImCBJ6NrouySCuWOsE4UYRVRBlYiyn4azhrgvCZdSstY569gwAMQQRaQsKwSUlFQU+zpySgTZOjylFEI0hsuiiCFJrmkMKKAxJkAgBAZJKU1mZ7WPEdC6orBoGQlZgAXYlOPhaFSUpau+tD9/9fX1OsV08F7we23EgbtBsbtlK4TOb9abGGIOhsQYFSICmWiYOQuUFbJaXfuK09laGdEYPnh+ZHF0LzvIuoT+qnz45pap51y0EBQSRwQNXW928bCV+3SHqNL6EAXYutKSQ7CEjEqqoJIvXkARlaQphCTadN5ba6xlw1RaUzrjLBfOlM46a8j0r6PEwJjzEMC5At0wFXY65uvttlZvIn0PvXLEEUccccQhjgT0EUccccT3irIwFunibDYbD4RFGABBg2iXJHrfhabr2rYOsRHpUAKkqDEaYmKTi8IklaKsXFWJqjUmG2gW5aAajJAIrNVyoMQimrZ1F9O2brZN2/mgO5Ww7iYnoMCMzjADSAxNU2+39Xqz6QTqtm1CNxhGBQjBEyEBAqpzhTFWVGOMKftZqoICUl9IKoaQUiLsi6WrSDb9jDEmSaDZdpOZjaqkGNu29a0H2ZGkv1Ma+oNM64cT7j/CyDz4/X3t8Hecvh6qWH/zJg8P8NANBPt829+wHX5kRx+1GnjwwT+BOQQ++BtVRLeb+vrN1dXrN48HT4rJcHxyxkz1oLh5+yp0vtuulqoj1fPnn1k7tmRSCCl0MYSubRfzqxD800//1LrS2GIwnm7X67Cdd81mGX3btpdPPxmMRl2MiowCt7e35fi0HI6rwSD6gZ93q8UKlS4vL54/f75ttj74rvOIyGw29XY6nkwmUyLumvpiUv35549e3TUvrxbb+E8yPA87YjcifxMh/GvxMNLwsX0++PA7BF8+/mUA8G6pzQcKaMy8JiEOB9Vnzx/9+x9/8cmjWdjeps6PJpPZyUm93d68fRubzWw2GQ1LjH6zuGu2m8l4eHH5qGvq1epmvblRaBEH2WmUUGPwV1dvjCsunjw5efJUjdvcvb69eb3dbkaT00ePn9hySKib9eLNixe3t3ef/+mfXTx+VoyGaPjr//I328Wb6P1wNLl4/Hz26AkKLm9u3r78Zn398uzR5WT25IY88LfwYQX0Hw4QwCAiashGrbvF9314PyAxWz9bwmk1OBmNhqWrnCkcOwOuIFfQYGDKkh2jdYYNIyESExEAASICOetK5xBRiQHBGJMjk0yZpFLDTIzZfRhAClcYQ4gQgxfV0jkmAtXWd0JkbSbPQVMUVVFBVUQEgRg6AM2PHhVJPhCSAqQcESVIKSKjNUYlJVFIIYYUY4pJBUiJ0ZAIJsCmk8aH2/nq5dvbr16+/dtffvXzr199/e1V04CPIHD/xxARUd+SiowIAKmPtiHeXxn3rYsIuCOgRfeP5cP++Rje56D1QDOdKcK+tB4hqmZBLLQJfAObpjHQ5EqSBcP5CD5/dvbDtf9hMo9OJwXqwJnKMIEws3EOJFmmwlnVCKCIUpZ2NBrGKFkLXZaVgpiOUhJJCXs9NxrrFBAgiAohWWtjSqDqrDPWsjGZZY4xFWWRaxVmA+iqGuRqeNKXjqCUIoAaa5AIFLzviMg6G1ovIoQooKK9vzSogkQkZDZeNWVSWQJqKl1BZABNVB4N+eTkNAkq0ia8kFVd+/CeNf/3ht+Z8FoBVIP36+UKmRBAkgQfoiQAJKTsgJap5H0S2756594HHQAyK90LCACJQFKUA+p5nzWiOwp7bwAOmF3Y+wKoCnhoEYZAAhIFGu9DSkjsrBlYLq1hUEIhUCZEApEUU/DRi2gS8W0InTKTNRytCZadNd6ZUFhnjbPWWWetMYadQSIkQlFUkeCDJAKl2CnyH3ao8YgjjjjiXyKOBPQRRxxxxPcH/clPvt5KM2NnTQrtZj5v2xpQJEryMfqoIkhoDDGkEJrCWVO4lJwCqKKyAWSwjqyzzhVlaZ01xiIBESNzTpRNN1c+Rh9jiLLs9MWr5WK56Xz6oFDWGTOpypPJqCpc27VN227rpgkpiibQrusANIkwkyCqSIyC2CaRPKXoOi+SQIGNybo2SSmlJJKnIhJjJCRXOFWVJCHGbP0pkiQlSVFE2rbJk5Z+/vN+rua7M8MPzdkQ79fSXVrt/aKPEnOIpKAPFZ27nfYTpY/hHdHoO8JU7TOk9Z56ODj+D/7+znf29PEDkRwe7mpPFO06VHfTur327l7heNA6CgcbHu5UH/x4cF7vkST75s0Kv/u13iMv93x7/jQfaUq+qe/evFrPTGnRlFU5PmFmn2Q1v/FtLZu5JdwaO5id22Iwu3helhWSWdxct9vt6u7KsHmknxXDCVnz5JNPF6+ir1eqMYZ2tb6rRrPp6bmx1c3V23q9RlMMh8PhaDgsn4HC7c3Ncrmwlp999nw8nTXbzWZ+MxwMz0/Pl+vlYrUqijKBNm3Llp5Oy3/1fPbzF6Mvr+o2Js0sD9C7TGUvPss9JL14uG9A7TWPD4tE3dNTDwXFB83+zvB4bzR+QBb5zoIDbvvXyV3f0UjfR4P0flDtroedyG1PrOHhIOgZBiCiT58++vc//uJHnz8qSGt0xXQ4Ppu124X4VkJXFOXZ+aUbDW5efPP225cphSePLn2zLgpG9ttm4WP4/AdfjIczUqjXi9ev3pjSXT59Nn30SAy8+uZn16++DG09Ozl59PhT58rY+na9uLu9ub1dfPZHf3r59NNqMu3qzdU//HR9c73e1KPpydNPnw+nJ6oyv3598/JFu9k8fvbcjWcyOefNJip+D5kY/+xQlajSiSbYGQv11ChALsCYtc8gFmlg7LQsHo3HF+PRyHJhwDAYC2QQCJCZjTPOEBMws2FRbrtIxNZa5ywIRJ8QwRaWjQkxiAoAbJs6PyRK54xhBWFDxlAKbY5lqkRU8E1DhCKSHRucszEEFc2lBUUkBM9MzCgp5RNpmibGSICGGRFDjAoKpMBoLBfWokguX+A7H6MgO3YDLkdmYDzIqo1/+4uf//TnX/30H766nrfLrd+2Xe195yGlw+AhEqCIJhUFBCDoCWXI10u+QerBPRHueboHBQ/kOzGfH3wOvrul7tjsHZFIOUgpABEgARBAAkgCr7ew+Hr5y5uf/81X1589vfiTT588OZtdTIfjqhhVZujYYHSMheW2HYxmATHbXxhATqpJ1RWFSmyarYqIguSzIirLISJKjN57UDA2s/RERNZYNib13hxSliUidl2X33yKwiGgSvI+qAgSdV2XUlRSRCWmylZEnAMSOc6dxb6SBBARIcaACMYZixSTNG2rIISa+dckCcCyihP88Rd/NJqdeSj+88+++er1tfxORNC/M3L51wIPyhzHGJumnkynzhY++BhC1jonwERkrAGEGJMKZJW6iKqIqIJoCjEnse2fA6qa09dSiL32GQGJ2RpABJEUo/YGb/kZAIg5B4GRFNLO/62vHoGCgIAJ1CfpYupiGhgWTTGKQDIMxhAzWiZDBtEAVAKyL2WSa11KSinFptlut0kl5VZXIWOMdcY63pnJW1MOeTjbkts2HbhR5OYnP/kffvKT//n776MjjjjiiP9mcSSgjzjiiCO+P7y4KD77Wfe3f63betOEOjTbGDtElZRSSKCKoKqAbJiQDDOiIaqqARCrogCDsWgdsWE21rAmCV1IKYokFUVNGr00dZIUVSOau/n25au3nW+AFeVdP1gEKCyPhuV4WFWl6zpvrS2LEq0tODtMk4CKJMMGECRJ9mo0pi/VVTinqoD9VF9EmMhYuy+PHmPMno8ikjAp4E53AwjIhG3b7soP7mqm/yPxkMJ7R1Kq++X3/Br2ImLNTiE7PQ/ubEP2AiC4n5zC4daH/zz42W8OD6VtO25uT8Heb/4xhfIhv7A7kHflmXrw+cP5c38I77DMO8ntPWe9P8r9Cntd3Uen4ogPTk73bDTuT+5DJPbuX6Q6Gg6n45FBWd1dW0vDk1PjnJhieHIRJaUUU9c2q2UMaezj9PJZORyDxsmZR8StuV0vl8vFLTGfPXo2OjnTEIfTmWpqmzqFTjcrLgblsCwHg6KsUtIYQ71ZMal1tqgGo9G4abbL1ZLeWDYGFbq6tmxG01nbdevNerPdVmUFgCppXNCfPJ7+my8+XbS/ul61QTRLut5pn3sv13s6NveWqAIRAYCK7kbXgfIUAUFF77vyoQ3xA4HkQaxADxb2A/43Myj4gd8+3E331hv7T/XgwHZcJRzEPna/EYCqPro4+fMffvbjLz57ejJIXV0NhqPptBqU3eZ2s5wPqsF4OuWyXN9cX795yQCnp+fTyRQwrdZ3m83SOHv+6HFRlYCw3awXdzcxdo+ePRmfTAHiZj5/8/pXzWZ5OpvNTk4FsK5rB1pv1m3TXT5+dnJ2WVSlb7Y3r7598dWXMfrxyezyydOT00swOL+9ml+/6pp1UdjBeFLNzrZoQttE739N4/1hQFWjSAKN790jD3pXAZQAHNKQzbQoCwXwXVQiUWBQQUkQEygEH2zpjHBakwsAACAASURBVGE2TNay3Vk8W8tF4QwTEiKAcZYtp770ABhrmJmQGgRCJAJiYEZjiImJKElCRGsMKoiI94EImTlXqyPqjYhSjES5tBqIpBRjiEGSoPYDmIjYGjIkSVKE2JKEAKpMlASBbFWOW6Hl3fqbv/vq1V3zZqVfv3zzzeurF6+vNp34iLvH0uEd7/6mulePvm9HsN/kQ0+1nsrW+wfIbwv88Be/t1peKZeBEwBBiABtgk2d7trtXRPeLNtvb7Yn4+HFZPD8YviD55efP7usrEViZy0jGU2GKZ+eMZYBoygiAqIrB2nnhgGU/RsQFNCwBYOAzjk2Jpee3D0lWBhZhBgR0VqTJIEqIoCKiABqrizJTKqUGzkXjTQsaAwSomCSuGvFvjussWSIDYcYRRMhkGFGtsaooKoqkDPODUqI7GwDko/8Dwb7Adk/D1JMTdOcn5/nsp+ZW94NXmTmnMTGhokMGYohxhAR+3rV2tftpBxiyFHJlCSpgPaPLkDIXiv3oe1d9GVX/PMwJL6PwewirQACGFV8ki6kjsEAIqPN8mQGJMj5CUzIhIAmB3gBNL/Q9XVHoNg7iYAiAucMgKQp+Qg+OQcGAmHXoEhIYGJ3Oi/a2ffeR0ccccQR/03jSEAfccQRR3x/6Ar4P/5s4rr5ar2Km7lFNJyzCxGwl/+ISJ53uaKQlIB4MJoY6yAroI1VY1VUk0gM7WbTbNax62LwKSREIUgIoghqDBaD1Xb99uYqiGcDKKgpi896DowAnDHDQTkcFGXhmGhQVSEpOWdcwdZklXJmnAEhpdQ2bYyRuS9nSCUi9emcouq9z0KnrIzZn7iIxhhiTKraW3NkpZZKSrf9VKfXPv9j9Ud5Irqr464IOQM5T3wyIQhMQNzz0IRZpaYizAYJZccB7ihCwpw6umOncb8X3DHTOyZ6v979wr379SGBmDNRD1lE6A8Hd6LT/U76L35XL4s7ae29umq39YOvfahoxQ8s0/yf7qR5OwJaZXdgkKtn7b/2QOXczzL3Etn+PA6/+b5Xdi2nvQQYJc1mJxeXF9Op3W7neJ2ShNHpKbJzw8k4JRRt1otmtQ1pjeysLZ21bNxocsbEhOhjbJtutbw1hq0lZlsMx2gcb9frzcKnsNmsRMGaYnZySmzapm22a5BYDgbO2tlsRoTL1fzt65eT8WgwHMYQQ1IArKqqaeumqT1TVY1iVMfw5Hz81z/69OvbTXxxt2yCGpPDE4cDEIH6DgYgwjxFxqx2VCViAFAVRHqgFwbIhpt9uc48FnajaTdD3zMGO58E1T5igvvl9JFyg3jfdfjwCx4wXzvF9QcZtF79pvtj2GuqezsfyZ8q7Eg4Zvrijz/7qx/94I+enHJqUgyjydRZ2zZNs9mmJJOTk9F05n37+ptf+baZnZzMTk/ZmuC7u7ubtguTk8vHj5+DQL1db1bLEMPZ+fn0/NxY2qxu59cvQ7sZDifj6YV1ZVNvJPpOpO3aYjh8+tmfVGUlsVvevL1586L17Wg4vHj05Oz8wjK1zWL++uvQNmVZVYPxYHrmXLlZbdv5dbtZfR9m9P+sUIAgkkDl8KIHgPubb3ZNVQNQIFbMI2MgdG1q1WI0YAwEQ8agYWgbsJYKx4bZMltjHBvDLBoJwRreR/2QkQyxMfnuO55MqrI01kbfiURjGDQBSFUVzCSiIomIiqLQJHpfnzZHPJEN447mAhVEsJZj9J1vrbWEJEl824FqOagMO+tsTD7G0KUUOk9A5WAo5NANYTBbzTc/+/bmf/pf//f/8vO339yBACSEhCBAivRgSPxjH1D/fLh/cPVMtB5EVpPWa3+zvvnFixsDMK3sF8+n/+6vvkhcTCpzOi7OyFgylhkYUwwiiTNpqBBjBAQ2LkonIkxo2BBi6zsRQSRVob7OIBITIaYYY0zEpAAiKQZFQshB+JhQNVc7BIDsHA3QFzxIkrLrF7MpnAMAEem6DjRHsjk/gV1p2RgkCqGNIRBCPnhLNgEm1KhM7Irh9NXr21dvb95c3a63jRxW29y12O83diM2xljXtTG2KMusN8/m7PnTHDUxbKyxxlgiatu2BWBmJWUiACBEa22MMee9wS4SmRXTfahqtztjzH4FQACQFKLGpO/66t9HbgBAARKAT9KEWKKyEFpEAGYUgAQCiqyShexMBIAogghEmPeYwxjWMBujAkxsTRFCbH3XdJuu62KSyhXkXEKwjA5sBJwuPve8+F13xRFHHHHEEYc4EtBHHHHEEd8fbqfg1FsypS1aUzAREsaUlJAMgytcWRZFhSBk0JZOQRCUmUFEQ/RN7X3nvfdt57su+o4AGIkQLYJhyBnVTLRqmhTj2ellNfKmGPrIXbcnkB6oZq01ZVk6VxCzqIaUkkrhLGYK4ICWytXqiqJwznnvjTGGOaUEAEhYuCJPSPKabEyuqu6cI6JMQKtqLp7el7IhQtC6rolWv2Wu6kPF2I5+xVz2CgkRgTKvl+skZYoPc/l33PHKBP1vzIyI2TcEEPoaO6nnYQ+55T31B5lX3tPPO900AgAB6o5TfigVpv3h7b4IAA7Yxqw46tOzD0+v33e/C0Tq14T99kh7Mkl3H+meKt8xwj0Z3a+X/xbojyOT95rZxHwO90T7Q2rykMg8NILsVbM7Yvr+BGFHVecfKVxcnj9+8uT0kjav55vVLWI0BqrZpbHlcHJm2VhTeP+KAVNXb27fWuby5NyWIwUMMQ5DALiL3i/u3kpoTy4eF6PT6eyi9K1/9auu3qxW89B2s5Pzk9MLRNJ01zb1du1j8Kdn5+V4IirberVZL6rSnpxeAPB8vtisN9aZyXiEpN4HJhISQJwU5Y8+m/336+QGV282AYzLQY53tcy7ESEquKOoRUVVCDmr+6DXism+6YiIiFOMudl3Vct2F2sOGanuR8KOfc5aNt0P/T4lek9a768UPThC/JBU8z4QofuqVAC59BNCNu0WkZ1UcH/O+0BDfzagKpJDNbPp6K//4ou/+NNPTga8XryZzSaF0dCu5/NF2K5OZtNyOEopLe7ubm5uLs/OxpOpcUUUfze/qeu6Gp2cnjwv3aTZLjbLRds21XD05PknWJX1cr66eVOv7qaj0fT0mXOV75p2uwCIzdZbNzy7fDq9fATer+ev5zevttv5aDZ+/Pjp2eWFs6Zd3928/nm3uB2MToaTi3IwHYxP/XbdzG82N2+a5Z2KHDLs8IeFPIQSHJrH90EMgOxdpDmyRKCEOLCmMgjRIyqqAiMIgoCKgqAiCKhGAtKsdRTQBAJAAMLGsCEmIkaEfE/Gno9kMoSSYhcCMxkiiYFQmVFTjAIiQsSomoJXUVQw1qhqTElEkBCSVlVJRL7r2NpsG+2YbOEIiYBAKbogSdgaBEjBS/SoaoGKwcQUw2I4e7Wov/zm9u++/M9fvZx/+2Z1fbuYbyFmmbBCtmVQSAi/q2JlD3Mdvj88uGmrAoAAKEIT0y9er263f/+ffvrtbIg/+OTix//qB589Ob88HQ2JY2gltCRKxhoyXFZIBKrRR5VUGpsDug4QjWVjYooqkrwnayTFputkZ/WgoCmJsQaRcjljSZJ8rlQsucBdMsl7n0SYGQBQCZU0ihefyxd7760xzhgiBhER6UDQBwUM3idJiAoISUMLXUjURawD1qndvlz9n//v3/8/f//V16/nmyZK379/AOzzw0iJYoxxW9eiUpiicC7FGFPS+whELhtpAFBUUZWInLV9kWiAnLtjjckEdKakVTWmiIiGWRFENaWdczRz1iNTzuvRJEgRY0y/IbMkAbQ+rDY1FTYabEkNRmugKI1zXDgzKApr2DAZA8awYUcEihBECZRAfeoSocliezYqagCGFgfFSGGEiIV1XJTqHAxO7uruxaLxYcXB/W464ogjjjjiiA/jSEAfccQRR3x/YEoR4oC5KAqbBuwssokhAhmyzphcOKVQSQoSVUWipNAkTylijKFrQtf6rk0hRB+8bw0zGovMubg8KjKboiwSczTF4OSc5z4K+gghHYhZcW/xCUzsrMvEcdfT24E7rxCSSvbf6BXQkEkBAgDvPaek1ua5YvZ3RqIYYyagHWCeH6aU8uyxz5812WBQrbWSUgw+r/OeN+5vxAMGGoiIGAkz55zTgMkwM/eMBxPlOonM+UPCvDoZw9hzv5CTOpmMAqSYp+RA1Euhd7tT3RF4e455p3feGTPoftku6XRHEmfuNtPDB8arfYmeQ6np7tz2vbb7srwb3SXaAuxFtf3h7fiFg+RuPRDS4v6zHSmcaeLdJFx7In4/R71v6XuFOPQWDffHivfGJzsy8+DAH1LYKcxOTy4fPzo5xyItm+Wbrl7dvpVzOyhmJbkCZDwQeFK45e1tV9f1Zi3w+sQWxWjMzo1mp4jEgMu7G9+2axB2duJGpXFlWUya85frZeo8CUbfGcaLi1OJIfi2aZvsn2EMucINhkPv6xCDAFjjAOnV27eX52eD4QAQr66u5/PFbHYigJ1vZ6PqLz+7WNRer5taC1sUuUrTvd5cFRSIKWeL59EFmYAWzTGDewJ6d93scgJIkvSRA8QDTVnfHfeBIN2rjHd9upNMP+ilh54xDyIPh33Uc8+7Mb0bgaB9oCN3noioiO4EzvsO34+4/eaZPXKG//VffvHXf/aDZ2dDjOuu256ffooo2/U61GtVHU+mTHR78/bbF9+cnp6dnp3ZvtZZ+vLLXz598vTJpz8oB9P14q5e37VdbUs3OpmidbLdXL/8drm6G4xGT55+Ajhou9Bu69VyDiDGjc4fPz27eBKa1qCu5rddvS5LWw2n548eVVVZrxfffv3lP/x///Gv/vJfu8FJMZidnj+CGDfL5fzmej2/i94f3Ij+0Nhn6K97uLc60gfXeE5GwWy+QTQ0PC7sqLAVk0NwDM4AWzAGrSFr0DBYQ85Q6axhYsPO9PdbBHXOlmW5qw5A+ywLYjbWFK4AgBhDVZaGOcaOUJmBmHY5AHsFLBCSc05EYkr7kEtZVUzMxmQtZJZaI4EmIWBDNmXhpkbVpALGOEACZJ94uY7zt2/+/uXib795+9Off/X6er1cR8n+yAD9NQg7N4Nf60f0e4iHTCuSgiYVAuiStBt/t7n9+s3tqIBXN8ubpf/B87PPn559+uRk5LAyaBgYBDBK6q3tk08pRB+zNbT05l0phRBUBJl922Zps2qWv2NKEmLIj2NRTSGmGAGAmZm5bTsRYeaYEgBYa/NYyPbfCBBjTCmJiDUcmAlRVZJIzH7cu7Gzq+4AotQEWLd6tWyvVt3bVfibn3315avrrYegBGhA4+4p/Pt+1T84/iSp67oYghaFNUYVQoxEtHudSETEhiWp9AYb2QVaEYEQQVFJVDS7rChxrgCqogoaFTIBLSnbXiCASvb37ulrAfnN99Ec008KUQDIEGfXdwkhJuhCohBNCDF79hhjjGFrjOlF8moQLAKiGCJlAUPISqb38zHO5ldBayxbi64w4wG78vWy7pIi/uF7Lh1xxBFH/IvCkYA+4ogjjvgeQWrJusKVrqiKCQ+G5AoIAsaCK0AhhRh8iKq+69rtqmub4BuJgREsI6mgCkqqigLLIgSXUso6ZVBhRWNNWVXj8WRMVsqhvXwK38y3ddfFXDSQ+hpJO00sATISo1HB4GNdN23Tbbd142MSSZKA8+wi7QnoPMtXkaxjstamlLquy0YcvRSTyLmy67rNZuOcy/RDzqstiiLPG4ui8L7brFZ1XXdd94+f9e24CrKcWWXiXCaH2DISE5ksO86EIO4U0dnJgZldT6OryaIfBEJWUULJzPbOvjL7VkOWKYuqqOxJxh2VvCNZes5Qe8eJHdkN8CGK+YCcFdF7enBHMPdUzC6p9d4M4dB2Y88mwuGCe510z4Yj7ghGANADUgX3fGROdM2lgwBQD4wX9pwF4oGG7h1HkUPsU2zv6WwAAAlKSMh2eHZasV9gXN9d+bZdXr1iTeVwQuyqyclwMomKPr5pt9uwlvj6V+OT88nJaTUcIFOMUZS2q3lTrxdff3np0dhicnY6HE3Hs4tutZSund/dxJTOLx4Px2NBxMWi2Wzu5jeD0chae3p6LgLbur6+mY/GcXYy7dpNSCGmYjCYPX5Uze9uB8UgCQRfp83ioqAfPhluo/7iqqWytNbtxcA9pZzEWpsJaO7jHyQi2XlDVUVSDkOA7FTFWeCMiGbHfeB+RN1zw6AgOxnyPTd9KM9HoF7D3o/P+8gCHmjZdW82jYC6H3Wa2fD+g/shl6MZe+OezJof7rcfvdJvKyKMcHE6+Q//7i/++OkEutv1djmbnbY+WWopdY60Gk0RsF4vQrOeDsrLiwtmZNR2u7y6fg1E48nMQOrWV6Fdz2/fTk9ms8snxWjaNtvl1VXbbMtiOBqdeU9tu7i5vq63a2OsKDx69sfD2XkCBoNf/t1PY7slLkbl6Onzz0pXxHZ7d/X67vb26fMfcnU+Pv+kGs+SpsX1t69fv6hDKCdnw9kScQmQ9jGb78w83svMv9v6/zzQXSW6Axxcv6ioQAAMMDR8XpUnVTEp3dBZS2hRmRIbMAatY8NoGIaVqwpXWMvMxpA1xpgsee7Ta4xhY9hai4QK2nWeDRdFYYwB0BD8eDQqnAvBgyZCJQZjjDEmhCAiALm0oTHG5gJpxlkAiDHlO/MQyYcuRm8M58HYtR6QnCvEOvS+aYMCENliMCDjEvDN9eqnv3jxv/zHv/npi823cx+yxB8h9apnINzZHH0H+uz3EweUOpKCiopq7/hECBE1tLD5evHLb5anI/jTT87+w7//ix/90fNPH59ZtBhTCm3wPnOSKCohbJuNpkgI5WioBD6EEBIilVVZ13XnO2ssACSRGMV3vutaEUVEa23Xddm/azCoyrJazJdd5/NT0zC7oiAiVQ0hSEqgICnlDQlVU/K+FZEE2nZeVcmYsiyJTEoiCoIkZJeNXC/af/j6zS9fLX51XW9EWwXNuVhIIhEVCKivcfeHAhWNIbZt65wjpBRj27TGGkCUXMiR0BiTkqYkElOOzqcUc9pB/9Kyez/Jb33ElGISkRxK110wff+IF5HeyAshu7J8rEm1ryugCkrMRVmOx5NZaSsSCU0MTUytxNTG0DaSC6PkdzFEMMyWjWMqDBeWnDXKBhkgEljo3/gUVRU1PxpFVFDFMpSlxZSIRNP30w9HHHHEEUf0OBLQRxxxxBHfE/QnP/mHDW7GOBgNq2GJTePrZdqoRAkpBVFQjSl5H0USAlhjJLYgsSxtirH1nWF21jg3yO/ytqwMICIVRZEzJjGLzZhACJT8sqkX2+2qhSSskHJu/I6TQgABKKvq9PSEmTofWu8FlJh6zpQZGQgAjGGinFkpIoCYpwEAsK1rAOgrEKqEEPI8xPuoqsyclUpZBC0im80mU1fee0kpp1TnYlM7HemvxY7/fGi/iwogMQkqomCiSEKIlBiJEGImxol2tBkiExk2AIqAzHxAwGTSOGvucOfhQZyLZB3QuJmGzpQ27HTQSPS+5QX2phsPBdRwYIzwgLDaC5bhfk97mfVOAa2gh6aVO27xcMteBftQWd4Taniwn71Zx65hAVXvD+J+N/ea7vuv03fJtv1X9xLt+0TvwyYGCX67rVerdUgnw+F0cnqpKW7Xq3qzUJXpaRpOT40rgGh0egYIy9ur9XIZlncKag0Zcyoi05PzrFWPMcQk9Wp+8+ZFklgMR2dnlyuFdYxN08SYAHA8OysHw1FKMYTFcumDn05ng+Hw8tHT6+vrTb1p6toZnp2eLhbzzseytONx6Zuu2TaiADGFtj45mz4a4UkRHXR3N7dgTB7YACCSdZPETKqaYiSmnN2OO+eL3CKEtGs7zKYVvanKbgXsQxq7zrvXJ/dqvp0JTBarImC2kiHqbRX6EIPce7Qc6EnvJX4HA3IX9rgPL+SRtpeAIj5grmGfLoC9kHsnkU4xTobVJ4/PPrsYD9lTbLng07NzNq6t176tnbHT2QkANNuNpjCbDInJOPbder64Xixunz15PplMU+hWy9um2brCDUeTsnDJN/P5dVNvAMkVA+ayaf3127cp+kE1KMrBcDwdDqfGFBLj8ub61ddfjUbVeDyaTMeD4bDeru+uXi3nN1U1nJ6cD6ePXDVOSdbLu6s3rzrvi8FkOKuK6ipfX4fDHN4FfmT5v3TswyXv3RVw/4MBLMKQ6LR0F6PBwHBlqLRkUQ2BIbaWnGNrM90Mw0FZFc4aJkImNIaKsigKp6DWmaqq2PB9BgmCG5RZ5ZqjL1VRkWVgLFxJvdWFIhEhMjIDEHO+WIAtqqKqLUpVjdIiWyQUUTTOGmssEyGAoHGSJAAwkePSFoaNQ3ZN1C9f3/ztL7/5+y+vfvHi9uur9d02tEkEe555fxns7tC9Zvvg2ti15Ic6H9+5P/7u8dvucXdDxnxrAtyXR1BA2o8KBVVFURXQoJpqCC/Xi//t7//vv3vx/HLyw8+eXkyrScEVowFRibHzEjyKgCZAdF2Iktq2TaLMXFRlCCGllIMK3gcmI6opBlXN5ScRyBoHCF0XutarqrEmc6AqKjGF1MUYcZfflHO2YoxF4Ywxogkw20lYVSBCTRpjiIpUDDvlL19df/Vq+au327tNPa/DOkEA0pwLplGVsM8Z+kMLOKiIxNg27aCqhoPh0q2orq0xWQSdaxIiADESadqZSBk0KgqiWRSdjTj6zK3dkx2xD7gfjsJ82RDR7gmlhIQAxKwpakqQa2sQiqTDMDwAxNA19TqNsud7sihlYYgGxIqoIpGZjbG7ELyiKiFZw6gafNIEkaTDvr6oscZYZsPElMc5MyIbMHa0bpIdd77RXTj4iCOOOOKI7w1HAvqII4444nvCL0/sF78M/9ePC0AKMaRm630XY1QBH3znPSIqaBKQlNgYNxgyChsaDkofgoAYY1xRVoNBSgKgxhgFROLBYMBMqqKIklLnvQpECc1mefPm9ub6NnXhY/PUsixPT0+ttXXr27YloqIoASmbYiDfGyioqjHGey8i1trMIHTeE1FZ/v/svdm2JMeVprcHM3P3mM+QI0CQBMlisVhd3VqrL6QLPYQupOcpvYIeQ7rThZbGpbVaQ1VXi8UuNgcUSRAgkMjMM8UcPpnZ3rowd4/IBFjFVjehAhibi3kSJ8MnMwt3t2//9u9cVWOMaf0rAMYQmTnLsmTKAQBJB52cPZnJe4+E1lpQlc5AEP+Rud8XgNo+FCRKQn0gaSoNJILECAIJQGN3bsmHNFDsiB6CIUaiBMTTdCtB6rTEMzHowSAZAJg4lfFJkm/oaxV2qtHTs0Skbpo2qI6PZLaDyv0WHTPuG6ETrvafSt3QI18FxTfaC3slEvY7ehNAD44Nxx2f2P4ebTKoswQ9uYZO3jSccHe2esLQ+/2eUuo34Lee0C8ADc3+sN/uNnVdTUc8mV8CCDDvVqv9bpM+OprNTTbKx1MiAoI2xqY6lPu1ZSJQtNlkdolAMQhEydyhLg+ru1c+tFdP3728etRWh7quQoit95vNBo0bT2fj6cTHUN6Uh0NpjcnzfL5YeB+8b+umOpQ0m8+zfBSCNk27mC3ms9ntzY33wVhjGQtLVyPzZMKLLH52t/VoiRmAADTGiDgUzkpJDFRI1jRINHikaIJsqp0BecoKDXy4V4T17PfYf50i/guIf6IyRNh3dK+Z7v6XVP3dWE393g0Z6juqO9oxv9Ihqk5JjZ2qWvqhdSSw2uHnDkIbovmk+N57Ty4KpFA6xmKymExnZVlXdY2Ik/m8mM2366UPgYlc7tBA5av75e12sxqPx8+fPGeh7W5f7g9IePnkeTEaq/d1ud2u7phHo+nc2jx4vz/s66aaz2aLiyvrRqPxhDKnodmvli9/86tyv7m8nM8Xi8m4EF/fvf7s7vY1MV9dP5ldPB1NZsG3u916tbw9VNV4OjeTx+O2Ypt9ro2/JtHB1GFInWSZkro9OW8YgBxx5swid/Mic6C5wdwggzKBI8wsZ85al2yAcZLnzhkENYaMYTaUOc4cK4K11lpma5BJVTHl9LirFxdjRGRrDRMZZmMYhhtN+iIQIJF1DmAgTkqIZKyqshW2FhHFe2OYTKeLBFAk40No29ZYZ9mogI+4r8OHn61+8stP/5+f/fKDjx9er8paQJL3cbo5Yt9Mw21Yezr1hbz5KxjdDQffyKAMa2SGi9T+piAACBgClOvmZv1q9Alcz/MXd7v3rmdP59k7l5NFYTOC0FQSfKpCgIQRMMRYV03K0caYNMWoEkKIEiJZTv0Yo6RHJFubboLee++9yxwRJbeNtKypaTXGmDnHhokovWwoqMscMwFKotKukBhVowQf2iBBcNfq7a76xW+Xv3yx/O1dGQA9YABSIAVAiKpDAuJrGKoqMbR1HWMcTyZ5ljMlFwuDiN0anCgCyADCnJ4haXUMSP+2IsniBlNtgyGdSX3+FU8e+idY+fitIgWNIYZuWRfi8ZVINZWbgBB805QhNBJRKTJjZsgZZgNIoGqY2VibCg7g8PqBmFh5Wm8ECJJeRKNIwssxRhVRYcNIXqiJ7LCA2Hq25mva7ec4xznO8U83zgD6HOc4xzm+pGhz/J/fH49i87DaHaCJ29tErKy1CmCMYUbrrHOZb72IElHmcmNsVuSFwngyQURrXZ4Xvb8DtN7HmNxko8To27at67qsAJ0Xsyr1Nx998usPPy6r6lT8NJwSAoyK4uLiYjQab/dlVVUuK4pJRmR8jF4CG9Le1M8YMxqNdrtdXdcJQANAqvgyGo1CCCGEPM+ttQB4OByIOMuSy2domsaYtIl2Ff9iTB7Qm81aJIK8WXjv3yvSdSXxcV/irzcdlpOJtSIgETrnkOiUzhIzEolKKkuYNKoDYB2ASD9fSmW6kJAiKgKQUneQXtvcHx0wnRecTreOM7TkLt1TSxDRGEKqhTjA5J5od/YbicIkqoinXEQ7EnjknF0D0OX7tQAAIABJREFUnM4Iuw1hcGropnDDlLB3NOl9NTS1YQ8/ezEvQLfM9ghMjxudcPZUIq+n7Sf/E1/XkxDati1DbrNiNOEnaJwA71YP++0q+DqGdvHoXTCW8/FooY+Y71+/aPb73eqeYphfXMt4lhWj+eUjQq42y9DUVbkNoUGA+XRijBnPF8Zmh/U6BtlsVsg0X1zMLy6qumr2+7qqyv1+NJ2PxqN8lzVN2dRN5erZ/HK33R4Oh9l4PB6PnOWmKQFgOps1tS8In02zZxP+UOuqiYJGcehVGcZIT3h08FQZrJo7E4seQA89k9jQ6ajudgh964H2+zgKmrtmT7tSAAA5UUx3Q6XzxxmqX0qfoYDTrE/XlSd7j5KWPcReHni8iaStuqvT4wU+vrp45/HV977xZMQBondFPpsvrDWH8tCGsJjPLp88hszVNw0xG+OiqsvNxx999Pr1Z+Ms+977385tvnlYHTYHJHv96On06XuxPtS7u2q3jk1VXF5P549i65f3r/fbzXQ2uXj0eLG4ZpM3be0clcu7u09/ffP608lk8vjpk4vFIrTVbnV78/ITD7xYPJpcPpssHqHKZnnzcPNpVR3G04vLx+9CcZFt7pB+H0XcVwxaDGSVoCus94X3WgQwABnAiGgxyqeZy1EzQ5lhx4gKBsEyOqKMOTPc4WZjGKFt69yNitwhE4DUTcVMqlE0WHFsDRI5k1lrgsQQBVRTPVtrrTVMCCFG37bBB2eTw0YQ1aR4zPMcEXfbHQAa52KMRDQajYwxCZPazBrLTVOFEBXUWENoJQgXYzZ5VbW/efHy737x0f/6f37w8euHvW9XdSwFhsX3A4j9//wI+grFPyiafkMZ3/ttoQJE0ADgWy2XzWb3278v6Onc/PPvvfv9bz759rPrzFiNbWwaJjTGGGdVNc+yGEVUu+wXISJaM7HW9uVMsWkaiZENIyISp3chEQFQQiRmQ8xEotq0bQghy7Okri3LUkRd5gBUNLLt8spExvtYHpp84gLwrpafffDx337w6Yev98tDaAA8ogApUlqBkp7R2uUgvpapJwXVtDRtNpvleU7ECUBTn2IUkuSXwb2TenrPGB4E/WsNxBjTEyJ548CQ0x4O9oUAWpOSPYYQJXqRqCrpcTa86SiAqEaRIFER2BgCQVUVCV6Q1BhGBY2REC2zZWOMAYW6btiycy7LMmuYkWIqkGgMMgKBAkQRBc2LTBHa4IvxKNjM4g4V3nn98MfxvT/HOc5xjn8qcQbQ5zjHOc7xJcVqxlccD1EikIBRzp2z1pgoQoiWyDpjjGEm6xABiJCYmJmNUQCRKCGKSH3YxxCCD963SZ3bbGOUIDGG4CWKKqIlIUvOtRF2+8qHqEnJ2gPCQXfJhp1zyV3DGEPMlPTDSRQnkhTA2i+3Z2bnHHFX1S/vZZPE5MhBr+WcTmfpX6iX2xhjEnpOUugYY9vUhxjSks7fqwWHTyF8EQNCSmSVOseDbrFu/weCMhMbY61JhY86LtMbIBBaROCkEtUOriWPjnQAUenI71GY3J+adhYVBHDUy2EPeTXV9dOeeqfjooggoJzw4eTxe5QWY0eEe26QTBsGyDmooXsueFJnMmFrJe1b7ESSfAKgT6eLPaCE4bwHmgzD+Olm7KfybRwO2P/XMNgGPeHQhx3+yjM7GuXRt5tdOZuM87yYGmts5ly2vHm5eng47EoyxeTimp1z+ZiIIIaVvK52u81qicg8muaTeTEaMVBbVaPJGCCUVf36xSci+vTd9x49etzW7U3U9f1961sCYKT55aNnT59vHu6aw6GqDnc3Ny7PJtNJlLDebB4els+fjxaLxXa9/vCjD9958jQfFwIxaXzvbu/Q2OuR/cHzxad3+93Letd4Aey0z8ksWQRQmahv26E5hobtrUukp8hD63WjoOfZnUP0G/g+CZl7r5ded3ZULh/hc6caRQQUpFMTGDjt3ONg6ZMQR5F7XyZx2OgIoE/G9rClYf7mO8/++Z99573rGTTLSGqzsctHVVVKbIEQrEPD6uvoa1AxxpDh9X73tz/5yfXV1Z9849vO5r5q2qpmdpOLxez5txBIlap9tV3v5vOr8fQSldar1c2rV3nuHj96Np4ufNTal9PLOdW7ze2rzephMZ8+e/7O7GIeVTbr5c3L3zZ1M3/87uOn37i4fspgDtv1ZrWuy3oynj159t54dlkF1taHpvmq4eXfK7C/z37u4rD/VyQABp04e5lnM+cKRgYxiIwCqghCiI4wZy6YHbNhIkSIARBza5gRQDDVAySDqMZQlrnk32ystc4xMwYgBFUt8twaE2OQoIoIKs4aZ21ap2/zLMmljTE2eT2PCtHkDUUIoBBS6k4ErQEmDaSKqSoCEtt8Ml9X8fXdy5/+/Ne//vjmw0/uf/Hp7epQR4T2TauFk9v4W41zvDPj25/9ygfiW7puHQB0fxcHPElVKEBUlACr0NYtbGtq5Ga199uy+e57zx5fXEGoNARUsc723sHpPgdMlJYNYXf76tytWu9VpAPQSMyMhAoQQqBk8QwI0Ll7BYnWWgCNMbrCqoJhTi8DAgKq6cM+qMlGkbL7Xf3r168+eLH69c1uU4dGNabqDDg8QrVPykKPWH9HcuarHRqCDyEws4J639YVpTZX7cpMqwIQpTc0SEU+UsqKGPun9um7wunqKThZTaHdKhnofyGggAqoGkIc3kBU+xztyUeDahniqqwcE+eZMoBBYiYQBCCyyfiNVUlANYYohJhZkzmXZQ6JDIMhIOeSUzT0JjoKBgltZoBA1FhngqWRVWH4L/77v/6DN/85znGOc5zjJM4A+hznOMc5vqTIc1APbIzLRg4CgIxHhbW2qipEtB0YBVFxycwSO8ATBBAUFWMIbV03VRmTaUBV5XmeZ66qqhhDMkskNi4r2DDZLM8nalzZStS35F3dJJO5m3I0Tdu0jSqIiATvQ7J01Qix81sUiRBDCJKcXmNUVVYFRBGpm7or8YcYYwTALMtjTFXvFXr/Dex8kikVFEqCmkEv/O/Dfd78KHaiXgRATNaEAACDh8bgkMHMzF0BeELojDWwI+DJR7uXPyv13s5pXWdakJwUU6cK1P4UetuC3j/hOKU94rvPEY5UEVCG4m8IAESpRbqd9cfqCKL0E7+kspXecaEnxX1j9nuDNyVvSZUMvRHDEVYewXg3UDq/BQQAoJ63D7Lb9Mn+EN3PIybvUgQKCqKqg7lozy05mVWoIIS2ripCZpNnRUHsgzS1917aurl/9dl+f5hdXBWTqUaczK4KN94uH7arh7I8yO2nk3Y/nl5Qlo8vL4hBkaOs2qa+f/3CWitBs3z85OlzJnq4udmt1igAiuPJeDQaBd9WdeVlM9KJdfl0fgHIy+Vyu1mOihEbNtbuD7vpdOqc2x8OVdNOppO6qTJo3l24f/knzx/KF/VdWQZAImYgICBVFUQ0zGllwonMOVUpVDwOk2PvDOMn9e1Q6++0cYfhQD2E7saX9AOABizcc2FK9SQHoARHnw3FXofYD+A3l1FrD93SlygpEzsX0BPh9unmzx9f/+m33/nOs4uZEwQzml6OZnMBqvZ3EOvReOyKoi7L3fI+HFYkGjFvQvujX/w0z+ffeP7+5fxxU5Zhtw0SxvOL2fVTZAtNediu6jrY4np+8axtZbd92CxXIDAdz0m53tfIPJoU5JuHm1erhwdEvH769NG77zjHu+XDZrUqq3h5/c1Hz741Hl02ZRPb+4fb27ZqJ9PHjx8/mc2vAKmttvVuGZvy982HfaUCYVC96+lvUx4rpe0MoEWdOHdZ5BPmDMGgGlRGAQVmtIyOOTOUG3ZdChIgRjZmVBRgEEEI0FpjrFWN1rnxuEBENibLCmJGBEIVIUUocoeAvqkVkIjYYO4yY0xVlgDgnLPOAWIMASQiwqjIQgwhBCZN+UtDykygQaMoEEJE1KSqDBEboA8/u/3bf/er/+1f/esXr/ebg1QA4eQejPD2X95snSOuxzeeOF8fQIkniP0t+oxdHvWN70J6eDQAPuqhlN0nq9W23pQHO55MLubT8ZRjixJsyjYzMzMSKfYvAAAhxhiCy7JUriLGmJ7LkJ4LRECoiL5tCTFzWVcfFTRKjBIBQURjjAXkAACqSAyIUYOKaBSJCozR4HYfXyzLn3z48pcv16+3HhkCQoR0VYPlV5cOPX43cKjd8LUK33rvPTFBWltQV0QJQKuqxhihK5PM6UGjyX9Du/Vq0MnSj3f+YVvVN54IJwnLFIKaxo2ml7237j7dVgAK4BWqqOuyzohzYLUIyghgCA0jxXR+gN0DMqoKM43GRWbZMkYJElQYrckME1PK5QMioSE2TAaQCYmMwUAwsVSpAsDP/uzP4Oc//wP3wDnOcY5znKOLM4A+xznOcY4vK1DtnI1kF/N5gcFCYQwTc3GxgBjBh7ZtYgiqEiF4kaqu6qpu2iZ4b63JrAm+adu6retxXjhj8jy3lpEwLzJrJ3mRp0J7CsT53PMklNQG2pUapJ9In2geDXMxyo0zIYayqdeb9aub1+PZHNms1tukXBYQAVHpFkuKSAJqIspMho0CqEiaRhIRMXvvJYpzDpFUIcYoEpNtNAB676011toQosQQg49RiFgldlz194xTnp5kcR3qO6Jg7UXHAtKLYSBKjLGGAUYz4SAbVjXMaExajEv9elQYxGLY8bsBKSa43fla6FGT2glSoRMFJe6LPRY86l2xVwefMBHtf3cCfTsuqUcFEQ4yZD3Rsh1VriecGDrLDezo9HD2J7BywNrHvWqHIFDxZNdvYPeTIx0x6XBgVFRUUhw0sulSFMAAdmUtQ7SEIYSm9dYVJivy6WLmA7Ot99vYNvvVAyM6a61zNh9r5gEoiqzXD9Xqrg1NCHE8ezSZz4u8YGNUVdZ3KrBbLdsmTueXV48eXVxdtlXpqwpBtquHzBnnrM2zsqlb38KhnJqsKCaIXJZlbEONtTF2PB1vl8vReFSMRl50fXtjGFWCZXM5dn/yfPTJfdOE5d0hKJssywhRNYbgEcA5F2MMUURichNX0WRTQ0iIlHi0Hv1YO2k0IopIypswE/T8FwcJNA6e0p1ZRLejjhcPpQJhyL4k3fqp2P04AKDbMPlEp/8Wkf7cALtj4aDcRsBUX/GEogMCWmu+//5733vv6ZN5nhs0pshHY2Lb1NVut3HWjMZjQtysHh4++620bVGMG9/ertbbzeG73/ve1eLKV22zLyFKMZmN5xdk3GGzjftVbJtiNFbKfOT7+7vV/V3w7XQ6n00XICgilojEr+/ul7e3wYfpbHZ1dZVZrrar9f1tU1cXl08WV89mi0dAvN+udqtXTVXmWT6dXk6mlzYvlvc3u/WqKXfeNzD4qH+Novvqv3WHPRkPDJARzqybWlcwW9Tc8CR3ziZspXnmMssZonVsLLNJIlbICpcXWVHkAqKoxrHLncscIlprUo04a5x1WYghxJjZjA0xMyjEGA0xqBrCzGbOGCIKzCEG39RMKKK73RYArTXj0diHtm5qNtw07W6/m0+nhulQHrI8y/IsqAAZtJnJZ3e363/943/713/78U9/+fJmXVYePFFQjelelC4ZYTDNGdoBTrse5eTXfxTxD1xqp2TtPoeIUKm+2jfVr5eV/7vPbl79ix9+71vPHj2+mFCMBJFA0ksBEiGCiAYfJUZJxXuJVSWhZ0RsmibGmGUZCqaKpkLovVcRAGRj2BCItm2rCqnWpIrGGGPUILGq69aHKMLsKq+rvf+/f/z3P/nVZx/flHeHtlGQCAqg1D9eUTqDb9Svef8iAmHdNt77UVEUeW6d0zfeKzSliJBITmTNqiqhe6/rILUCm5QqECIePnm6qz6XmuIkKSpJTI2qktb+DNumW1JyY4+qIWobQuNb9BJAdhAdkzNEBM6ZIrejLMsMGyLnLDPGKHVTty1EiQCCpKbi3LlxMUpvO4zGAVlOxwdVsURsaJobafW//su//E//6q/OAPoc5zjHOb60OAPoc5zjHOf4kgJR/b4tCuMIMLRRKt9EUY2IGoJ479s2eTJYw6paN21dt94HYgNgka1jts7lWV64zLIRFbbMlgEhFZYhIgAERcpHIrasD1XjfS9JOaUqyY9iNBo550SlqqqyqlrvnQ8MlKYiIQYyTECSLAVEowoKKIJEUVUVQKKELFUhhKghJtBV1w2zYeYQfAhxUFU2TRujE9EQgkpUCcnwcTit3wF+3hSgnZDX4d/T5EcBIHbelaSdU6EhBiIAjSKA3YxLQUWJhJLAGQAp7RcFIRl4iB6rtOFRHnYExHBs2eFET3Fyr32GAXMMuunBhxkBj6rlt691MH4G6G0Tuosd5nm/s+nw+EP1pHZhOvtuVqg67L37AzvnDMJBCffmDr+QPp/S7uEyOlStvbKbeowKqSgeAKh0tsgxhiiBjTEumyyucpfXo/H2/vaw21a7jXN2srhwo0KIbDGaXFwdmqo5bHarVWgV1D599i4VE0QKvvW+sYhNG3frB+/bLLez6ezi8qKpMt+22+2mGOXFeOLyPGt9eSgP5YGNcy4bF+PZbN7WTQgeIBR5jkRVXbO1xhljTFMdENRlNsuL53n+g280q4P3UDbgsjwHVInBGIMAzMysRkXTFSKqqGETTCQkxNT4ojqoyDsAnTI6CRan+fOJU3TX0IOsv9swWXWoDF18YuRMiD18lh61nFh+95/vRlL62MCgu36io0QwbdVV5UxXkqSLSI+vL37wnXe//exilltCKYqxcy627WG3rZt6Mr22zjZNtX64a/Yby6b1fr1v7u/Xzx+/+97Tdy34/fpBvJ/OLybzS5PlbVPtlvf75e3l9cV0tggRt7v9er2sqsNkPL68emTdSAGtc1nGMTT3r19s1qsiL66ursfjot6tH16/2m+2mRs9fv7uaHyBzOXhsFst18vVbDKezRaT6cwYbKr9/d2r7b5qgtdeV/61C+xJa3/bOH6fFQEsQEE0z7NZno1zm2HMLWeWrSFmQIQss7kzOVPmrHU2KViZyWaOrYVEd0BF0LdRtXUui6h12YiUCMjGhhiiRJdZYwwRt20jUYjIECLiVpWZiLFX32NTNxLj/rAHACYu9ztVFY3EHGIM3jd15RX2+21dG1fk6HIPcAjy2e2rX/zm1Y9+8uHf/+bu1d3OAwiiIg552C6LdyLAHFrpC9vu6wopPydxxs/97phj6jXSCr2EWAF2Xmrfxk8fdk27rOEvvu9/+N13ni/GY8Msvls5ESMkXhyiRgXR2AYJUUH7NUjoWx9jZGRiAtUQAgAIdyk6VVWIIQbfeAA0ZEFVQmzbNooG1SjqA9YB6+g/u9384qNXP/7gk9+8XG1qqBUEMOpQWW+4eH3rAj/3l69ovPWAVlBsmqbxrXM2L/I8c433yR2qsx9TMEzEHGNMb4uEqJrMdLpHPCEppr6QPm89yKIhrbTpBdGYHnCqChIhFeDV40PnzaVhJ28MAipoiBwbZ9gpWFBDxjIxqcQQvbaoEKVlIlRnjbFEhGzYMAImVzIVVSTiEIiQiVQEJWoIFk2XOgUkgMwYp/7PfvazF++++yX2zjnOcY5z/LHHGUCf4xznOMeXFVGRiCWE8hDaVVOum7Zu29Z7LzG54wETG7bJixmAQMG5bDq7yLLCOpNnbFhBokYBERHlzFBmADV43zYNKhIQEwGS9+Fhud6XJRKA9OIlPDofM+FoVGRZpgpN04QQnMuI2Bh7cXHRNI33viiKZOaYXDjathVQ0c6CAwAS9U5TxBBC2/pUlb6qKmNMKkLILETYUy3NMpdlmfcUg/dtVBWJsbcG+EIC/dZvBoCCgwlEwnaACSN36LOj8SKYOSDsaCuiNSbpTKPEhDrSAQwzivoYOdFnRcHBFlkBOpNpBBBRBCCkjsp1Rh54ojHtWXFv/gyQzKkBOrOQk2TAm/6/p4X7jr6L+oZv7yDEPiGTetp42BP6YYNhhz1FOIqf32hmVERCwJTMeFPN1LPz0w1SC2F/8p/rstNFu9CLx5Om3hlr2XlfEyOCSvQSGRFsVjBZUGyrWqLU9eHu5kXdHK5BkVkJs+n0Mb67vqH1/d22WlrKrhdXbAs7nkyvnkiU0FTWtbv9rjqsl/dZkefT+YwNL+/vmrZ8WN4uFEbT+WJx2bS+Ksv1aklI19eP5/OrKis362VdV0z49PHTzW6z2qzzUfHoyfWr39YIwOxcVjyZzf+0kbttvfN6swdnrYJGBO6kYUCsjCaNfBUVFCa2tiP1nWoZNFm+nK5oTt0ioidq+m5iDydK8kG4L4KoStqPxk6QNrADSKRbUHsbjw4oYK+sPo6HAUCngpb9DtNaZqJjVxISMhIRAYpq4cz3v/utP/32829cz0YOfIxZPsqd2aw25WZlXZ6PxzG0+81DvVtNi2wymd+sy33VzuZX/8mf/wVKvd/et/Xa2mJ+/YyzkW8O1XZZbh422/Xlk0fGmrYu23pHFC4fLS4vH02nl+WhKZzJx7m1UO232926Df5qcj27mEdpb28+W97d5vn46snTycWVCB62q+Xt7Wp5rwjj6WJ+scjyzLeH9e3L1e3Lg9gW2I5Gb7uTfl3iKF/t/3v4QaAZ0sSYiyKfjfJpZiyFnNEgMoFJoJnJGna5s84Ya5jRWOusRcSoWPuYaFX0PmoEhMlEmCnGcNhv27YlIlFBgjzPk+61qioEGBVFnjtVXa83AGCtyfPcOWeMAQCRGGNI49IH75zN8hyYiNlaK0F865uqrhqltnVTs6rl49v9//i//9VPPnhxt4q+93ru0dhwYxwybyctAfA2fNR/7K9fq8DTW7ge04/d06p7DgGkQqdRO9VqAHi9k2W5+cVnm0+Xh23r//N/9v478yJTRUCJsakaSKldBRAF0fpQKYBisr0CgG7hRgveGCaitvYisV/8gZ5bSYUvQkTgSAICvvVNVUVRJbbFCBQaH16uD3/7y9f/y//1d5saDgF8/+4zQNHuSgdP79/d41/NOE2Gd3+qSt3WrW/YUJ67oshDlCjSpd4VQNUYNswBNFmeMKKi6YtfAAD0pt4gcnwpkihpHY52tQa77H43liRICGQMIKOigvTjK712DUnx/v1HARQzY8aZmxZ5rj43WOQZo6qGtq5EBETKqo4xqEZjyFqb5y7LncusMcyETKBIAbCOwkqsajAGVQox19w6aw2HoEBITBgJAEZw94ftk3Oc4xznOMdJnAH0Oc5xjnN8SUGIpOqY27aUugreGzZmZIL3WZZleR5DRAAmci5DJB8CACNZ4iypiTX6IIKglEoxGajrujm0yB2OCm1o6qbal3a02NT4qw8/uXlYtgKib0+ssIOLaNgUo3y+WJSN39YByRIZNJxlmfc+1Y6yxgCAqoYYm7aNEo2xqp3zhjEmy/IQQowhhJiclMfjcZJJMrMqZJmTLpSZrTXOud12e3vzeiBr0CuY/9FAJEAC6I2foYe62JsV9HQ2TYWMTRWyME16mBhSmZ3OALrjekxHE4/jFOtk3q0hyYM0HUnoaKmRGN7RgOPIdxOAVuhl1YkddhudSoeP2rNTjnsEyCcfAkgXc+J7gf2v07UMKmcYxNMDhR70S58rLNSfiQCQyNFSpKc2gIlo48mZdKpdOMqohxZ7a2rfOZGDgLJ6icJImTEakVXFe19WVtG4XADQmPFiYUhH4+L+9uVyede0LZObLBbZeMzOOWNi42Mr1WFf7XbL29d505q8yIuRe/bO6v6m3K+BIPhmu3z4xvN3nMlilmVFYfK8bvx2v2ebT6fzd56/e2eMr9uqrF6/fv346VM2pi6r6nAo9+Xi6dyQqZpaAUaT8aMnj9er9aGq1R6uRsXjEX33yexm295tV1UJSKggHQFOalDVEAR67V1Hd/vGGobZ6XrkgUQncH2SgOidZZLKC5KiGY69m5IuiGmUQVI+Q6pq2eV++iMqIgpKp2FG6qTP/Q5TloCIurXwfe1N1WMtRUDAgEykCnnmri5m/+KH33l+kZPft1Hy8VhBD+uHeruyhudPnkwurjb3r1naxWSUISBziLJYLL753jcLhsN+F+tyPBo9fv4eT2dt2ey3283yfr9bfef9bznLq4e7+7v7+4eH8XT89NnT6fTCe2KjWZ4ziK8Oh/0Kol/MJ7PFTCTevvjk9auXeTa6vH56cf0YC7f87PXm9q7cbo0xj58/u7y4YJRquzzsVpvlze3rz7ybRxnneYFfLwCN0K86AOhAYicW7P6VATKky+n08WR8NR2NCAgjI6hGHyICg2BAbZt6vxeVYC1neTYqcmM4jV+m9I0kplTFFlPpMmuNYbLWGWMQIUhQTfd/22UuATLrnLOIMJ+DMWk/aSkPhBAQbZ47xFSGrkUEZrZ5JqBt66NIUACTTxcLyosPP7v70c8/++t/9+nHr+8f9tK8WWnwzRvoQN+/Vn39HxxvtIae/OYLWD2AQrrfQQvgI1QKP/3NXVX5w2r1F+8//e47jxwTxuirqkOSoiraFS7AISHWHUNEyroCACbWlJeW5BBNzlnftk1dB+8J2LJLyzOYuY3qFeUQbzeHj29WP/347sNXy2UNtYAHjEA6vF0cL+ePqtO7Kw8xHg4lM89mM0XyPgwLqRDROcfEISQ0LQBASIj8+d2l1zhmFtUYIvaFHNMTv3t+iQJiqnrAzAAkPmpKJkmIb/tE93sG8KptiD4EiQFIUUFiQAJGmozG3bKf9KJIkJ5dyXZOJOU5UgVgNsZY2/Rvg93rbiq4nec5M6HN922oyYQf7tzD+A/aAec4xznOcY7TOAPoc5zjHOf4koIQkQiYBVHJ2GJsmYlQVbIsy/Nc03s/kWFGgBBiqtceBQgiqsRQqwYAQEFQUISyPlRNRUxkDJGpy7oqq/JQFWI3JXz64tVytYn6xkwSjkontMY4Z411gIjEWZYpMCAjk2FWkaF4YBJsMnV16p1zIjHxLGNs4gtEmGSGnhU0AAAgAElEQVRriGitBQBVtdYiYp7ng+OtiCKCtY6YBiV1r8T5PduyY7iAyQy5n2Fgh98G5W4nFNUk2+m2FU2l8ZSos0KAjiF3qC+5P8NQra+HOJ3VgWp/HOyIKw0nf2TBOuDdTnh9Kl4dhNC9E8cJYT6huwOR7uXLcGKecLSi7q+0PzwOTs9Jl9R7Rw9a6t5wQ08PfKKfBu3L0506Pp/6Ww+cfNhKe4frAZr3Z3O8roF+K4a2bQ777XatY27aVmPdQJ777UEAR7N5MZkImPzySgyNfBNU2qap9lvQiCgjM4sA4+nCsdutl9vVw+2rF5PqML28Hk1nJstG80XQkIdI5AzYh9vbfDxyeTGZXyhnVVXVZbVZrUD18ur66vJ6u97sdodmvy92++lsNp3NfFuX+93q/j7Lsqapd9ttPh7Nr64j4G63je1h8+Cnxfz9R/PX2/Cb2+2nDzvANCceciAA2rm+YG+XksTQiXsNxTFP275D/McO76Xux3HTtfbQcTpYuAz9nj6DoAI9fZYYZRDbD+kK7BZZq2qqMXiiUleNMUqMMUYY4PiQWklfQiLDdHE9//Pvvfu9p5MplxzLzObzcV6Xu/XdawSdX11PJpe75Wb58rNYbSdFkU8WZRPH43GWFyMr9eb1YbMkZ0eLR2Z6Cb5t9+v9eul9vH78pBjlTdvcvH7x8tXLyXT27vvvFzYvD03b6HQ6c5lFaMty+3D/CqC9fvLN2Xy2323vbm+dKxZX74wXzxTt/vbV7uGVhDhfzEeT2Xg+N9aW24f1/cv95gEgZgZH4zyEIjf8taNTA3QbngPHrzwDOKIRm2mWTfLMEZIGCT6gCApjKvSFSIqEABJD48UIAhJaZWZiJKI00pUJmA0ndw4iJrSGnWUkJIKoIqrMbIwxxmR5xkTOWgAAFeecdTY9OKSvK2CsmUwn6RcScwVFRJPZtMpeIqoBZ8eHaO5vDv/mZy/+5icf//iDl7WA13/gefIWRf3adfh/UHyeQb8VXyCjD/2wulkdyrKOvlpt96tt+fRiOs+t1SjBSwioimnBEWJUjZ0LkaZ0lyrUTQ0AzNzdsWJEgmQi7ds2tB4BDBrLLSIjGzI2gCkjPGz3v3px97OPXv3yxfLh0NQAsaPP9OY5//H1dZ/UDCHUdU1IeZHvD6Xvc8SEnSH7wJ2BkpCZBtXz53fJiStjel4dH0ZIKCICQkwArKLMBIARUCMiaEupFuQX7FUAIqAX9BFCVAFUTrUHEBGdNZxW3KAmBUJXlxkkSQWUEEEQU01gZuY3tPugIUb1bQQ1hjBK6zVYyHZTP/L/8Zv9HOc4xznO8TviDKDPcY5znONLilTLRdlQlpvMjjOjGknBWSMSJEaXGzYMyBA8qFiX+aoKTdWVFUMV34bgY4zeS/ASYwixFQlKCEiidNgfghdmx2RV493Darc/AMBb9Hmobp8XmcsyQFpvtg/LVXko2ThkAwGTBYfLshCCxJg8GY0xAoCE3rcxxhCCMUZVQ/DHGUgfaQaZcG0IIf2FmUNo27ZtmuawP8QYVbTXd35Op/2PRYK8p5C0x3GaxD2qAAJtCB1lJkQmxOQ2KGwMAsQQkTqapgIiwmx6mN1Rv/5nZ6YLb9hm9G7O2vNWTBeExzPqjCr0hMYeOXL/qV5bOvRT3x49OT6KZI9H7X8OOzwBlYN47UgM+yMerYfT/k+k2KnIfCeD6j8+/FQ4FjI7kTF9IdHuyGk/icWTbUi893VdlQcYjUliQFZyrq2afVmHKGSNLYqIbMaTOWJWFPvlw2Gz3qyaVA3JZEWWj4qsMMaotMuHe1iLMeSssaMJW5uNpiEq6kHbuF2vy6qcLBbj+cVkfpGNp6ubm/qw367XeTFyLhtPpj7Idrdbb9ZZ7qy10+mUQJtdSYhEZK2t63o6mY8nE99W281DW6lDHpvxk4l9PDa//u26AQRkOOlmRGQi7W3H04DqMjGnX8lhAAEMOrIUzGSS225vx6l9iHQ8v8s39B2UpOtdf6kqgIjGKOkrfNLnfeqnKzCYThL60+wAdAghAWg4WYUNRwCN49nknUeLP/v2k5ltKe4tyzjj3MD9zUPdVLPZfDSZSdDV7X172Bv1oJmwA47zWWYN+nJdHZbWcXFxVcwuY9C4X2/vXjWHQ5Zns+m8Kg/L1cNyeScS3nn33YvL63Kz3233EvnRkyeqfr15WN69aqr91eViNhk3Vbl+WALw9aPni6tnxhaH3WF9f9uWh/FkPr+4LCZzUG2qw8Pd6/X9DWi4fvToOhKPLpodaAxvJAS+JtFXZO2q6nW3FgJggIJplmU5E0ZfHypBMSionhEMkWc0hozhoshdZpCKLLPOWWYYFflkMsozZw0zECKwoTzPTYelkRmZO2U+W0YmQOx9Y3FUFFmWZ5k77A++bYxhay0zt7713guINdY5l+VZCB4iWGvJcLLyUISsKIKaVo2J5qc/+eD/+Dc/++t/+9tXq30ZO+b09erBf7rR+UEREEEUWNfxR79ev7jd/fKjF//ZD9//wXtPHs/H9b5syoOB5CrMRORDrOpmuL2ktVZZlllribiqqhACERNpK6GuqxiEyMzHk8xYRsjyQokPbYRi7D199NmrH398/5Nf39SiHiAACvavOXgyFv74xgQisTEi4tvWe68AhFTVdVXVqkpMTGyN8SEkhcEJdA5fyOtTDj69IyWbpu59qzscRolRxKghQBERIURE/YJdvbHbbvkbRmAv1ATMEKLSkVQIIApFBQwYBVGJmZkMc1qmZ51zxlhD3f2FuavcgekVEyKiD8G3tcuYnFFHIZoGgFr7H6Olz3GOc5zjHL9XnAH0Oc5xjnN8ScGISDwejZQYQxBFEBRUEfUh+rZp2lZEYgyxbUHVZlZDCG3TNhWqMkGPcQHAABIyWbIAbKwlY5DMYn4ByITGji4bLifTqcuyN88CB87FSLnLnLUiut1u1+t1WTbGRiQTkjmy6uFw6CSQneiXoBMw9Zro3iZwUNkM9Ln331AAIKJ08glYJ0lmXZUi8Q3q+vtFshY4XlD60as+EXtZcSJkSCIRRJMEvSMwqipCSojEzESJuaHAEZ4m8jiUjFNVSiWTgFIVnqMu9YhvMUlYeyHpCQTuW2lQOKueTIzxZPPTK+04YS+IHWSxR7ON7mPdNfeMciBoqZuGjTva2C+YPRkW0C/I7Vuvh8lfIJPWkwm9Qp88GFS7g2j8lIofUxMAYDmtzO1ETIhAhqw1oW7rqgoA5OzMEBjLxrmZHeWFJePbdrter5crFZ1fXmfzzDo3pmnUR3Xb+OpQ7dbWmhEhkSmKEQio17LdhRDa6AUBmCeL69l8Fps6tm1d1avlcr5YZHkxm0Hb+sNhv1nbIi+szWazi22AytfW2dmoKJuqrvbOmsyxxtg27Z63XND1iL79aPLhxWhZQ0Tu0h59X3RweGjkY4N3auLEkaErCHkyHIb0h0KMMYSo/ceG/x/zCtgvTU4rAAABYcDKHa8WORrGnAyjIW1w7LZj5iB96xmOF9Httlu4bfmdZ49+8J13v/P8gsIeVbJRUeS5tnW937h8NJ5fGOOq3WZ9f5NhKIrcuiKAIWtHBtUfdptVjOHq+dPi4jGya/e79e3L7eouy/LpaKQhbh6Wd7evY4hPnr7zznvvS5TD/uBDKEYjY3mzunv96pPd+nY6ck8ePyUNq7v7/XZ/9fidq8ffsG5UleV6+VAeSiIzmU0niykSHZb3q4f7h7vXbdPMLy7mj97R7EI4v6m3MXyxPO+rG10S683vLfb02QEWbGZ55ghYoiElVCS1bB2TY86csdZYa7LcZZkxBq0zzhlr2TqTOTsqcmcYAIxhY4yxnExikMAwWcvGWiSKEpEQmFTBWOOsA1BFiKrGmbSIPqoigMtyl2WiEmM0hm1mkYEiGWMQSQGC94BMNm8a+OT18m/+7hc//uDFzz+6vdmWVZCvW/99FUIBIDl9KYBCI3J/UHlZkr4oD/5f/uCb83x0URSkEUTSLc8JZEWRag8CgDE2y1yW5UTdywMAOGeRVCS2bcNkDFsCjCGEtjXFCG0elX79cvnzT+5+/Jubj282+6gRQAAFVDVpZRXgH2OfX+9QlRgUkh9GTOsPYtv6psH08qYwaAWEOT2gJUYAxC9SQCf/DGMVMX1pAyCkNXAqGkKQ9I6qCgAxJt9nJKV+HYN84RufQnpca+192fCeFT1AIBGbWwbmWjUziAaZ2FDSN6Oqtq1PBlMxiliOxpDhVJSQ0+OQuZNFOxdVfZtbyyYbgR19utxVLYDF//Yv/8v/6i//uz9oP5zjHOc4xzlSnAH0Oc5xjnN8GfGr/+G/ibElVMsUomiMEaLEqBJb1RC8Dy0AxhB827S+RYCiyEFFgm/rmlENs4IiEhOzyYgZAYiAGbMsY2PJWGMzQoPAkYuilCzPmT9/n8c0JSPELPk7o1Z1XVaHphUFBtKmbZiZmJNqJsRorSUi7/0pgE4Gf4lvpb80TZMmMDHGJGga6FcIIX0+KTq99977EIL0bg8AAG9h0d8Vqgr9Vj1IG4Td2iO0jplRpwcmIiRGwk43TZAQOQEyUZprJc/bJAGlPpAwhigipheihhAUYCiRBHDqp4F4wqbT73qtaQ+YOyx44oR49D7AE2SpR4Z4NAPuNzqx4Ojoob7RHqk1jkLsNxow/Xmiex4+2qF4GkoqHv/Ez+0hHavzcEgf63/Ty3jpDQuJDnIajMzGumwyWzBWYozJC84clE2Isd7thUgQHj17J3ofRQy7xfVjRFSg7XK5untARWOZZzN0xk7nj57T5vZFud2E0CrC4uoxkzXjmQETAxBy68vysIsxWpvNLy8uLi9D0y7vl4f9XhUvLq+K8WTqQ1ntl3e3RTGeTGd5kU8fXcJ2S4TOGVDxTQkRLeNsOn9olk3tp7nMM3w+4z9979EvXh8OHqn/xvV4WAdtcq8y7vTpCT+LKvRi5pOxMAwqAIXYAYKUTej+HDygsSfOqQ+JqUsTDCLnvsNw6K9Et6GX0vd1oJKF9GClPnx5hz30CZG0E13Mxt//9ns//M43niyKcrXKJ/NiOkeCar8qrJlePcpHs9a31f5+u3w1HbnF4tn44roKjlHBH/x+48sDTRf2+jlbF8p9Xe4+/eTDkXPz68tRZu/ubvabbX2orh8/ff9P/xnn0/WLT/br1Xh2+c43v6FNeXvzyerhJYFMp9cuG6/vbw67tcun777/AwBbblfrh7v9bkvEo9nMjcbIWFebV598sLy/F6XJ/Gp2/S6NrnNqvRByi/rFq86/0nGq/0xjINFnA1iwmVg7zVyOYlEtkWEwjJk1meHMcJFleWZdZq1l69hatpaN5Tx3yas5s8YaBhCXOWtt0jIiKiEaa7LMOpchYRtCWhGAhM5lWZ75tlVVILDOGkNN0xIxG+ecI0JACcETARtCskYNE0dRH0TBROHG029eLn/0s4/+p3/1o49e7e52MSBEBOnutX+Ebgv//0XKb/TjTBAqrzdtjM2DRl3MJz/45pPLxdyRoESQKAlSIid6aDi9F1jrDKjGGGMcE6G1BglVJXhPyIRU13XTtEgGXVGDvS+bn396+zcffPzBZ9t9G2NfRKJfogOpAGF6dukXgs+ve6iqRgFEjTF4b4zNrEXtiglqsnBGHBarpU1CCAjpWaanr1i9ALp7/VDV4H06SCq327YtABITQATQ9OIECoQGMa3P+YLFCdq/sUSVNsYm+MaDiUqCojEGEwwbUG85z0xmGSxhMuPQGIIIoGIMIkl8bcEqgiGEpMtnIgQizJ0DRE/MjC4vsunidtfsg59OXCy/wO36HOc4xznO8YeIM4A+xznOcY4vI7y2ll3T7OrVWkEQWjbcNHVZlofDAQCcc8VohMRE1lgiYpcXvm1AaXY5zp1xzhlniQ0iA1IMoS5Ll9tslCEBEgFybHyIERW8+qqt9+Wu9o0MKuG3jDgQCJUYjTNsGZmRgZ1F4rptRJUAnHOICN5nWUaIPgQRQaaiKJqmqet6oIpJJpnnGGMUka56obUAEEJIZh3pk3meO+dCCDF4773K6eT194YGA1ftoRoQd4JRBSIiToX+EInSwlJEJMNIpL0omI1hIh5cB3ppaF8ksCfIgGr01AEjWV0nPfhJk/ay68SQj3a6PX0+sVCAE7Cr6YQGWwOknkC+EXosNYeDUnpg052vRvrkCYAeJpCd8PktMW7/oYESD/rYtyeKb6UG3pxCHuFpB1cHmn08Veh05yIiMURjzHQ2LyZjE7VtmwgaEYyz4/F4V1Vt01S7w43/dDqb5XmugGTseHH5GIGYV7e3Dw+3aJRIs/GU2NqiKCbTtq6qsvQvP43eT+ePrRuNxhNis1mtbGXKclcdDjefvZiOp0RsrGVrEHG33yPb2Xw+Go1ms/lhv2+9r+raFRkZns7ndXmo9gcmaA67BnVcTB4/empN4WsffWuRvvNkjpPrrf/tJw9lJE6WmrFbIkDpwmOMacqfmkJEsOvuxIxxsITuyTAOg4NFRGNXxFMkSjdkEghOBjLDICbCY6riVPzej50+t9Kz5pNvVKpfeNqnKp1Raxo0iSb0I0C///63/vxP3nu8yMvdvURvspxdUZXb29evHj16PJlOyWXlvt5u7lXaKE7QEmfSeIdYlfu2qlw+unr+TRYNTX3YbW5efVIetlfz54hxv1tV5e7h4eHR42f/L3vvsS1ZcmWJHWFmV7h6MlRGJoAECiW6FrnYX9Ajfgc/gpxxsVePyY/g4pC9OOWgB6wm2bWqqlkCooCGSmQiMyJDPOnqChPncGD3uvuLTLCr0I1kJeA7Il685+8qNzO/12yfffZ58sGHZTULq/bNq5uT2ez8/DymsLp+HbrNtC4Xs8mji4vU+88/f1NU0ycffMjlZH27vL+/32w2zObyyRM2pijL1fLu049/8fknv3j25Omjx89ttUjkqpOztFynbZeyIcDvGk+lO+p5uFkCMKJRdYSLqlpUVW24AHSkhUVnjbXkGJyhkrm0VDlTV44ZidEYJBQDUBp0zrAhBNWU2CAjEKiCGGZrrXPWWsOOEZCYqkmVPYqMtUgIiEUxyfEpUNCUrA3GFM4WiJA9Y4qiAEgpeecYiVLU3oe+j2Trpk+v3y7/9f/+l//ub3/6dr3pggQAARAAIADJuff6BRr6yEv/ZvgS0vDXASHXh1NVXXv45O2av/czS7Coiycn9aSsnWVVFUUFDCEw82w2kzSEqIkpp0mllFJKzAQKvg/b9WazXoUoxpXzi7N1xF+8uPqzv/7hjz69/fSmaUISgMNpweA5M17479pn+h+B3AQYU9quN4vFSVlWVV33IcSYQIGQnDWtSBy9/of9EAkxyVAkIz+jAFCzvlyzqFoRQEVD17Mxw1MFiZBAZOhjACRkw0wIkiR42U3UHoQEVEEFERCIyTqLEIOk1HRbUAY1hKUxpbOF48KZwhpXOGMJ0ZKx6CyiKqMwpzwVFI2SCMEqEwERJbYAEHqvBKhEdiYJYwJ/48DFL7TbEUccccQRvxUcCegjjjjiiK8CCtrKlkAJUUUQ1ZCiNVzXhbVorS1KZy0CakyCiIZdUcQUJQWjyRJba4iypwQnEUVyzqlK2zQpxSQSk6KC96FZt256dne/evX61Wq9+nVLL0Z01hFhTLGsyvl8bvtkXElkiqKAMRs/pRRCKMqSiCQlH4OoZnK5KIqdY2Beeuzsg4l4pwF1rphOpznTNheH2XFgMf6ahMz/T2CW6MIBs065DGO+BiUmw5yP/FDLTMikIzdqjCEkVaGRkssa1exveMi44qjyhSwYHRVAAHt69VCYjLoTRe8OsV/aHaqSVVWVUA/4xAOt8H70ZBfpnUvG/sJg77cxaJQe7DjuPf58eEGjpnqvkNT9PjBS2wfk8o6/+rWCsnwERNTdV9gn/4+yb2FE41w1mbqyNlGQyRa2rCqr3PdBmU1VXTx92m8b3/Vsna1qkEhFUczm8xBiDHdXb7ablTU0SeImc1dWfVXX84WCtpttu1pV5ZTYItuiqmi9cUWNSIabvmuvX7+spvOidI+ePFmvNmxj8P1muZxM6ouLR86VXduqyna7KetqUlUgqd9u2razhoLvWm2Qiul8fudvfdeTMefTmVTltx7NVm242oQ06Na/IBzedcNB0w1U86iPfte8ZdCx78cGEDGqEu7G2k4yfyCh33e4Hg4ChVxsUFVFEFEOzgLjkXB/0eMIzQcjxN1xDdNsWv/Jd56/dz7BsNn6+6ePLiaTGQD5kJCZrW2aRlrfbO5Xy9tJXV88flJO5l3XY9/54LfbLZvy9NGTYjLzfd+s7u+vX2/v7p89eTaZTGL068369u5menZx8fyb87PLJHp7c7NYnC/Ozpwpmtu3v/zZD5H8+fni4vwMFT/79IVPfHLyuJqfpnazub/ZbjauKE/PTucnJyqhb9b3N1dd2ywu33v64R+QYug7LpA0xnbjmyb1LYHu3uTvAg76d/dCjoMZpIp54uzEmprJAjjWwtAgcyYtmArLdVlUpSudIUJjqawcgAIKDU8Qa9gwEzM654w1AGCdySpmIkDKtwJlwqQqqqIJIogKWEekWd8qMVfr5AicUgRIQKKCqtGHjpAAMAb1Eba9vPrss5+/uP3RR2//5u8/fnG17PIdBmEYzQPZ/qWdeGSffxs4pPXHrA8AAfUKt23EV+vFTz7DFP/L7z5/enGysNYaskSEnJylXIjSakocQsyu913XpxB67421qtpsm7brQlKyRTLFKsAPPvrV3/7ss+9/9Ob12m/6JFnqvA+xHPgZ/Z53Oo6f+JS89973quCKYjKZDKH6HPhkzglqgKiqKUbI5kuHHyMEABDRXD8DAFRFYpSUVCVn4jDR8KyXYQZJYyVkQMz5ZKCoKvju/GF4QGq2y7DGAhaYZQuKoJawMGzZKEpIoJASeE6EqFHFp6iamMAYcm6YLFtD1nASytWzZdsgYEpRmYAj+phENaknD+H3e5AcccQRR3yFOBLQRxxxxBFfBUSFkIGwKKqUkBStwcqVRMzGQFGAdZAixKQhARMwgyVFkBTjeoMimjSGmGWuISZRNYbbZrNtViGG3ofeR1tUfR+ur25OHqX7Zff69ev1ev1wbQgwpKUCE1VlycjBh6IoZ/O59QJASMZam20BcbD5S9a5vFJpu84HDwCZfX7ITuKhXbL3vut6RCwKN5lM2rZNKTlXpJRC8Jm5lvSbeEADUhZc71LKicgYs1MxE5FhTikpwG6FNTbCKDQmyjYmKe5qr+GQX4qIRLDzSh5lzbtibQ+v5pCpzhUKc1mmA/Jvt82eMnwAQlIYy/Dseioz3YdGCrg3QRhtF3Zs5gMJOQKNR3qQlLz/TmT328x8ZmtOGLyAQUf/6Ads6Z4ZBX2XmIZ3toRRkJZp58P3ywYAURCRLaEzJMYaYy07KMsyqrqqnk5qo3B/v5T1htkUhUXrMPpyNjtXUQm+3d7f3qakC7JFPbFFrXMFwBRSu92sl3c1YFHPjauqSe0Rmdkai7BcL+9CSrOT87qeIXLXdZvVqtmsCWF2cro4OXXObTarvm2JKdvU1HW9Dj4lr6K999BsF4uzoiy9D6pakJ5Q+vajydv77e262bQhF2bKwyxLvd6p4Kews+Z48OLhkDgQiu018kMUJPukHFQmHBpac5AChtGRgyAKOjhOq4ikNHq/4C7KcNi/cDCeBw3hqK/OHyVAgMIVz5+ef+f9y0UJEBrDeHZ+XhVl6IMSTeZnggSSUoq+bWKIJycnJ2ePinLSbTZxu4p9R2zr+Xk1P1fVfru5e/N6fX9TWnsynycJTdNsm8aU5dMP/3BxdpkUNutN1/UXTz+oJnW3unn74ld316+ev//4ZDErXLG5b29u7s+ePF+cXGqSze11v1kywezk5OT8nFFvbm9vb992fVvP5vX8bH7x7Pb159vtemGM9ptmfRN6IUg7ifrvCg4Z6CHYkdlZJqqMrQxXhgsii2oZnSVr2Fo2CNaQs1wVriycNYSEzpq6KgFUJObbGhM756y1xGCNNYaJ0RhjrFFJIkmTKOb0fEkiSQQ9Z6ejnF6TUuq7TlJkttYGpi4ET6zWokiughmSqAhowqBm2aa/+v5P/uL7n/w/f/95CxAAEmSr38P3e8RXBjz4O46u8ckQQbdBY0jf+9mrdrMxhiMAMM+qorLMTNk5KOtnmThhAoEUUte0TdP0fW+cS6Lr1VoViR2Xk6WXl9d3f/69n/zdz1++XIEHkCGShgCDDxfunnp4MEv4PQUioYqKSAih73sANMxVVWUpgIjEmErDMLovqWqSpArZ8C0/E3L2TVa2i+iwr0oKQSXt07jyI0bSbhzobgKUHyJsRFKea3xpryiAEiCzZSqZKucIgREsoWNiwhi8SFLQEGMSQNIkSB6SRCJlQ4WzlokQqrIonKWYC32waoeAjJCsSeRi1/VRQhK0CeV30HnpiCOOOOKfJo4E9BFHHHHEVwEVRAZXuPr8XHwPfkMokAuyiITNJsSEKpqSphSCTxIBJaYYQ9QIjGQMGwYAkRSDjypqnWm7TdtvgTAKxCgpJGT36PJxMVvYdfbBI0MypFEi6EgJEoBBrMvCWasCXd83bdt5IbaAads0ogKjLbCqQtciIjN3fe+9BwBrrTH76uGjucLobsE8UtjkvReRvu+zE3RKyXsfQui6XkR+EwL6i82rGmMkJkRQARp9DyAvnHaUbxpWRYjITKKiCr3vmdiOizERtSaMOtCRgAbYWx2rAABC9jsYVKc7nnaQoI5+HDsD53yAnc3COxc//n/YSWN9uL0F8wGlu+Ozd8rZnQp2vNS9TceoZh5/cygQPNSNwah8hdHp8YBS3l0kjOzmntIfOW0VGDXUumczxwuAkUxHjACd99uuUyDNSduKKpKJWmssEYr3zBxD6NpWU1icnRTTCSK5oijPz6yB15/9qlmv9f6O2YGodZJM8DwAACAASURBVCUZS2RA4Pbq7f3yNoLOEZF5NputFUJHhtmgrtb3XbtBZkKqyikCdE3T9P16vUFj5ouTsqr6rm3bpm87VCitLYsi1fVm7RVZQX3oet9WdR2j+tBL9CTdsxk9ndHHFN9sOyWCfUvl0UIHvbzvQxxfxQPj7HG/wWdzCAPsNlXdredxGJb7YMfBMMjdMh6ORgYgV5oaY0WZM9BxaO130/2PY+RFIyRVYaK6mHz3m++9d1rX2KDF+ellPZ1CTCKeDReLc0mxdrZrGg2ddfVscVFWEwLSEJr1PZOdnz6anl4gmdhstve3y/tblfT06WOVuN2u1tsGuHj6jQ8uP/h2avv7q6vtelXXk2Jaq8T7u7dXVy+qyj66OK+Kqtl29/frspg+fvxeVZTb5Wp5e6sq8/lifnJClrfXb371yS+2283i7Ozy8XumnCqabedbHxYg3erON2tBC3joy/51x04JvE9cyC8gKIGW1kyrsrLGIZAmNsAGmdEwWSJDaA1bY6JITMkWVlS8j9ttayyzISYCoJRkvd4iqDHMTEwECCJRRIwlZkKiJFFR2XBOjgGmTEAPTgsh0N52nEBJISEKskhKkq3OlRCMofL17eZnn17939/75D+8vFsBCIACMrKASP4JAHR/e/2C/vvL2uiI/zgOH1jvaGLzXzrccl+hAVAAAuhNBz953Xb//me3TZ8An5zMFmVRMIfeS0qEXJaFtTbEEGNKMcYY+943bYvsgYjYuXLCRX3fhh/88sWf/fWPPnp1/3YLIcfxdqVU93fcg4vdhfkedPbvGyWtItL3fjJRYmq7brPd6r70gCLzYcnBMdiJY+FlEBFAMGxyONmM8yUe1NWSa3tkcnmcb8JuQgK5OK4KqvQovkvvRM4BsjQaQPOnWZGAQDVFJrQEVpFFSMGZ4bKsyeUICVEBlSm7UYGkhKBM1PZ+2zX5ySuqudwIITrniqqzva6S7aI6YT3eCY444ogjviocCegjjjjiiK8CKUkMhkrpvJe+U+8JksQokhAxxZhSBFUERdGua2L0CFkxBoRWkSVET1ElSPSSFBUkEGgqmMkaIANkFK1xVTGZdcmmeBujatq7Ax9OsYnQGlMUBSA2bbdebzabbVJSjJklzVbOOHrEeu9V1RiTGWQiSikheh1knsP2uV5ZFn6qakqSf5sLGIpI13UAICLe+xD8b8g+jyzwnh0F1KSqMhJ2/ECXPEijBiFnZqSjUF4q9X3PRGG071DVECLhnn/bqeuyvvuBe+/ogLDTkeb3CzDmIo8SUwRAOtjjAAcsiQ4+zqNwePd+R+J44KB1t8weV4q7g43+IvsXYC+b1j29uf8lHNp6jEUPdW/HATul9F7KjSPLvuPZs+nE4W67M+2XueNxU4ibbdN0HtikqIbIEMUQYu9VNfuhhCQhxCAppCDbVeO3z59/ULABJtCkMn/y/L23L19sl6u7N5+3m+a97/xhUVdkSgAWgtur15vlDYD2IV4+eq+qphIhtNHaYrE4WW1Xm/Vdimkxl3o615PTmGS1XtEKU/BVVVrL0cfkBaJ4BFSxlqbz8+12kzSQhbvVzXz2eLY4Cb5dr+66zX0Jxftz88H55OXtthdEolFcDpDZeQAAlSEYsI9YHAyD8QN3EMQYRtYhAT1EUWAsgol6OFr2fQRjpGD4Q0SIOgzQ/RB5ENt4OCp3g3MUUKsmkbpwzx+f//M/+dZZhYVSNTk/e/q4T+LXdxACcQluXhjDYd0ur9b3t5P55fz0sSG7ur25ev15u1o/e/6N6eLMFVUMfb9ZXb9+mSSdXl7Mz86uXn28Xt8HcGePnj7/zp8CFW/evLp+feWc+fDDJ3Fzd3/35v7qV4D+G994f1JPt8vtm6v7toc/+eP/wp2cNKvV8vpt23WLk9Ozy0dlWW7urj/++Y8///SXj9774On73zx79Ozu5rZr26b3iVidffXmc2NtEmr64JP8Rrekf6rQHQe9710CKIgm1k3L0jERCKhKUkFMkYRAUIUwgvSavFcf2CdPiMTQeiRGw+QK66x13qQkmlIOkDChcxYQAMRaYwwTs2hCAmOtqCgoCeXsirQjL3eewRpFFECIlQFiikkA0SIVqmbbwyef3f31Dz755Yvbm00fhnezl9/u3u9B+OXwLnbEfwp+HZm/a/yDJ8g+wokKkBBagas2dS+XbF8h0J9888n7l6eX02nfBt91wfvJpC7LMsbofQghIGJKMfgUJACzq2Z9L9v1+ucv3v71Tz75/i9fr3po057nPiCY94GWg2vW/WsHl/r7gYFcFZHgPTO5osgTsBjiftJiGBBhTFUaQthAB08hQMJkUjZxStmsQySXvJWUX+MhvWaMUxONcyXGJKKShih1nl89fGYhACGqqCSJMSVEIQIaKmYzAYGCKoEiAhEgKRHQUE0areFcJVpSREBjbBSfJCHikD9EwwTPGnZF6cqy8KaRDh4ErY444ogjjvjt4khAH3HEEUd8FYgxAPqmhbevXybfQ/KOIcWU7fMMDZ7FTGiIYpKYhFGZrXPWmlIVUopt30bfauyddWyMSqondT2pkNmVVVFNFBhsgdXkxau7tml9F0OQlEYR3MEc2xA5Z6wrYpJl09zeL1frtSsmve+QaDabZc3yLsd/u92mlKy1mVxmZu9D3/ciiYistZmA3rGHAJCLCI0MNQ3V51Ky1hpjvPcppt+sMUctC+zfFAIgqhIggY65oOPyRkeqNjtQp5QUVBNG5lxGfbgOouFIGndi1CxxzjwiQZZIpy9ImYeFzUAH7shr3VOue73qAXG775NxpTzQ2aM3wv79jQT0OwTzjtgdm2akLkfeGXcuGA+dHwaOE/dHPrzkvap6XLPvKOzMfeN4LcNRDjd44AEBgPuLHI4MSigxJhEVUQLwPqBKUbGkcH97c7/d1icnJ48f67Ypy6KqCzamaZvr12+mde1KpwhKbnZ6CYrX8Pnt9Y1PCi8+rWanZVm4erowLCmt7+82y6Wxdd82Vb1gNluE0C4BcD5bdN437TYEOQewRbk4mYvGrmu7dquni+lk+vTJkxhT6Lu22fq+M84+e+8D48qm2/ShWW9WrohuNnFc274Jt96wvHcy/ePnZ6+X/rO7TtkgYQ7JAAyjEgZjk/0Q3Q+jUSQOo0p99/Jhn4/k/j4EMmr8dBTLj6PmYHzCzosDFEAAD/XPuo8v7Aeb7uTzu9hI/moIL89m3/3m06fzklIDGlBd8nGzXZvQQYyRwHBt2Pzio1/4ze1kMp+fnFX1zG9X7Xalks6ePFs8esLO+H7bblbXLz+LoT87P5vU1cvPX65vb/uQLp4+fvrBh8rF5uqmXa9PT04uH53Hvvvklz/brN6C9heXF4+fPe3W7d3NOgW6fPLMnl02N9erm5uu611dn1xc2NKt1/efv/jk7dWrZ8+ev/+t75yfPVKF1PtmtcpG5G3TtF33/ofPfcDi1XrXX19z7MNnsBdBD2DECdmZLaZFYSWCRNEYUpKomhgkaDKJKBL0qCIRUdlwVRXWGVVJKaqmyaSuSuesscZKSk3TpBTZ8MliUU+qonAikhIAABIYNoUrsstQfohkCylmNsaoJM2PD4CkItE7x2VVbLddTMB2QmbSBbp/s/zo8/Xf/vjVPQAAEEJSVEA8MLl/QLT/xwXQR/xnxqHj0z7IiZgIe9DQyQ8/urq7WaUkzhSn07MoXdv2d7c3bTudTqcxxhBCCN4gI5Eytn2IIBOHb66Xv/jszV/84Kc/f7O6aiEgCI7c8t4Map+wNODIKw7RelRRH7y1djqdEPOBvZcioCYAAEkxP28QCZARNdtrAEAuk6FDAQEVFsildDWXxBXMrmO6I6DzvA+zdROxURFNUSSqpH11SIAHzzRATRCi9CF65EDojAINhaQBBESTCA5O1JgSIpJzlsgCABNZa7hw1hjnSmOZGWU4OtrCiWrwnghtOSlPL3DZ92+uhY83iSOOOOKIrw5HAvqII4444quAqIekhg1Ij+oBJCRAVECIMQJaREZCJUyEXE0Yp9YYayyzEQFrjbWcpFfpNfVsHTKDKhMZRFAhpJyuH0Pvfdc3Wx/63ktKkNmkPUMJuV6TRkmt9y4mBRKBmDTLmDWl1WqdLTUO+dOcMR1jyhmXMcYQBr1qXmoYYxBx563hnC3LMls/78iypJpClJQGavxL8A9ZMioMDPRInh4qmzQvhEYPg5z6CQoigKgECIQwmOwCorF23HUk80YKkHBP+eZGAFUV84D526kMYdiECIdl8Mi7jtrrnbD1oADguNtOpprX7iMBvZemZtI3v0I0mn7sSHaAbMQwEpe7UwxvbmQ392ut3fUMLTrwOPvd9hLZB1Sl7ltpJ/fOPMDAsQ4s+ANVNcDIcwIgoCZmS0QAGmOIfU9ikmHfN943qokIURNqSKE1RVXVM+eq7c3N2t9P5vNqPlckBa3nF6cJouJqtV4tb5HQ2TOwNVosp6fep67Zru9uCuessUzWOu7WkRCqqq4ns6ry26Zd3t9Wk0lRlWdni6u3fd+FZrNmgLKsEdFwnXs9xtT2gV1dACSRopopkSAyG1OUVT31vjsp6NuPZm+3aRNet8IKlBtUhn+6N7N40BWAiDsTzTwMkGgMfux7dmjokf4fXaLzan487DhqxpGzC4eMlMNIsj6I0xzosfe89ch5jxwEkuJiWn/7/ad/+uHzOasTrKvJpJpQStK1QAIgxuCkcpvVsmmawrjFyVld1aHrVnfXXbMpJ/Xl828W01nyrW+W7epuu75bzGcn06mA9k3bBzm7fHbx3jfcdNasV3dXb0qH80XtHDar29XyrcTu9Gxx+fgi9enq9XWz7SenT86ffQOi9E0bQyiryfzycTmdrVe3v/rlT9+8fDGdnV48fj6ZnErQZrVq7pch9CCBHQNAWVauLEUDaUQJvwtsBOawW+56QkAFGey8ASzy1NkSgYNHECQlYgQlAmZ21hbOgMRRVGiYEQmrqiyLwlgmBGK0dtAbls4x0enpnJmNNc5lcyYGVSQk4kw0k+EkSVTYWGOMYY4p5seKRBAAMgYIDWgKxAggWJUToULM5PPr9c8+efuXf/OzH3306h6gA4gI4wNAFWQXX33gqz6+eMRvAYdC43ew4xZRAYakmKSIyqCbBK824d99/7OuQ2vKs8oW09mCwDApQXZ8hhirac3WRAWsF2svL643P/z5ix/84sUnN+2dh3Cond1fDuqu3t07Y+Dda/y9GhVDnDmpdF0XY2TmSV13Xef7fpfihsxIQ+1G0cwz5zu/wMFDRQFAVDEH6/N0hUABokCeS6QhaJ8zfUQBVeCgCITu5qDDTzC+PkwboqQuhHXXYeIQaNNpabA0VBrjmCxRURiDTATGsDHEhNay4WwVoiAJECVqSKqBE2FWKyBiaJs8h0OiBOjXawPOICYA0t9QDHHEEUccccQ/FkcC+ogjjjjiqwABJNKqcnWBalxmohBUJbEnYwtbVKPeFgCI2RhXGjaEEEKyhorCiBaqHiUoM2ReNaQUAyRNmkKIkjSk5EU2m6ZpGx9FFQkhwbvrxKQaRKKIIrEtXFkXZTDWsZEsYSEyABBjzGyVMSa7aoQQRcRaw8zMtBNED8aygMzMHEWkLIuyLLNZh7WWAFUkxJhp3A473/df1lT/gMXh3qAgS3UAkAAQiBBIQYgImfOWlL9RFRFiIks7N+SBRB5JWBz5ix1RTA91zoSUSbudMPzB5Y5HQ8K9onhHvOal3s6zYk/n5ouhwxONklPdyYhh5AZh1DePRot7AnnQgj088zvtuue9d2fDcdvhhPtgxY7C1AeAcfk40szZhfiAVt21BBxw3/umQtAYClc44wAgBM+IxpisXjcGC7TWmBS8xD75zpa1q2rpQ7Buu1ohNa6aKKKyIUfV4uIMCMzb1f1dt7kvigKNUwUuJtUsimi3Wbabe2OLopoygbXG913woZoUJ4tKVe/u73vfTONsvlicnZ2sVsvY+2a7QUAyjgy7qkwqzbZbb5rFyUlVTVVEgfPFKxNbe3J+sby7ZWeflsUfPpl98urm83XqRDODvOPGhh4dXVSyEjm3iuxE4nu7jN2IeNCXQ8OO7pzvENCqo3f7rg93g+rAr2U3YPBLhsnDH3E39ICY33t88YfffPbB5cKkvnB2Op04a3zXsSYCNGVZVnVp8c3y1lg7X8zmp2eEtFnebldLQJyenFazhRL0fbO6u1rdXhvGxWzmmLbtVlIiU51ePpsuzkKM91dvUuzm5yeuxO3mZnn3ViUsTuZn5+eG3fXLz+9vl9OTy8XFYyazvV97H2xR1ovT6el526yu3ry4uXolmi6fvj+ZngOY7WqzWt77bWMtAwCDMhG6AkUgepTIqF9/dkp3YYoxqrAbAmqQCuZp4WpDTsUQGCLDyETWQGG5KorCsQgaxqIw1jAbQoS6rsqydM5k3hkRkBQRq8I5Z3KFTzaMCFmuiKiEw7MBCVWVhETVGJOTYDAgIlhrE4AIKgAZRsKIpJJE1BS1B7fq9Se/uv7LH3z0V3//y6t12wJGVNk/0IY3uy+O+u6z7uvfn/9EsX/QHHzdQ8eb/5h7A4rYKsROmxd3TOZkWv3RNx6/dzGbnp1iiioJhZJoUrFlwdaKQOjhZrv98cevf/jRq598drNU6BTk3VPvv/2S2NGBGvv3EeMTQEVGIzVblVVVlqDAg7IYslFa/pxKkpRSjuHryN7uni05g4fZQNYhg4pKDDHPBFKMOTdnmJwQShIdM7EUQFLmpcdrG+cF+bEFmKemGhWDohcVSKIaBUNMjsgxJU2FYWMQBVERDSSMoCgGVQgMqbICJo0SmYmGkDkBMhMRECAiJIl9T8YwAIc+5lniEUccccQRv30cCegjjjjiiK8CTOjInZ+dnM0dBAVRAJDRg8PY2hQ1SFJJqoJIyJZcDSlBjMaklELXdj5sRD2jxhhV1SKH3oe+3xFPfR8Ekcvybrm6W61SEiAkIonyztIsisYEbG1RVgb54vyRdRXSMAvH0cS567rsmJwrzKhqdtVgNiIppZRVcACQvaFTSsyLrJVmJmYOIQCAMQZGC4L829vbW5G0Wt7/Bo1JyMRmECdnmo4IkHD0caZsaTK8kUyhgogYy2z37xEBeKjJBnDAtRFxPmp+d0SDh+DOdpnGcj07TjivrwbKEGEsqrWvIPdAr6ogcOATMtLTu0UaAIxu0AAHPTfqUxEwF7AUHF/XL/AueddR1/zwEOM3h4cf9dYwash2BP2wkQ6V7mXcaU9z7gjog/McaGn3LOhwthj66XRWlSURiWhdlPV0ajn7krsUFRFjjMEHkcTWmLJsOj+ZLbpt023bjV2aspgtTmIisNXk9NIVVdds+67Zru8Bma0j5nIyQxCJbddukK2qFK6qZ7Om67r7ZUppcXpaVdW22d7f3fbtlhAuHj2yjOvlqu/8ersu65kBy8YVNfkAfd+KTMuyQpiJaNe2XVgbY1zpTk7OssbZKLw/pW+dV9fLu2UTFWjIQThoLARU0CFrYWi9vUhsGE6jD8o+wACwewkRQUQOFMrj3gdy5gNN6D5eA3hYolOVVA9MJw4uEkajFUDMCQeoMCndt7/x9NsfPJoXiqEtJ+eucBJ9u1kTASDXk5OqrJrNpt+sptPp4vyymEz79Xqzuo0pTWfz6fwsphB7v10v7+9uNsv799//RuGK2Hdd2yDAbHFezU416fbuZnl7/ejivJxUfbO6ffNivbyv6+ri8ePC2ru3V6/fXFtbnj97f7o4XV3dtD4Qmtl8Wi8WQeLt9av1/XVdusuLR2dnjxWdCHTtdrtaMtF0Ouv8JmrUJDFB6vrU9ZCiIfqa01VfIg3VPAABCaBgnjg7K4qJ5ZLBMliDjrFwXDhTWS5L4ywjOOu4LCwSECEzTiZVURREpCqiCUCZyVo2jo01zhoFFY2MlEN3NiudrQXVJBKCJ8TMPiMRiFpjmMkaKwgxQIjRILG1IOi9DykiuVUjP/7kzZ/9+x//xfc+2vrQAQZE2Rs9vBs6+fK74BG/dXwJ+wxweD9BAEgAohBBE8BHb27TX677+Mem+PAPvvnMQlLf+z44JHYGjAlIAfGTN2+//7OXf/X9j9+s2q2AB0iAY83Dg97+Yq9/rT/E/xkxsP8580WJ2FnrnLXWxhjHMCcq4s5QK08wDLEbtynLMnusEXOeBDDnitiqoElSjDG3eIxRhwg05Ky4vu9jCIgooklSiBhBJaUviNhBAQQ0qiKbcjIpDVUGSqOkiVIEiSGG5MU3agid4aKwzhpjiUiJ1BZcFrYqbGGtYUaglJJhdtYCgiJUZU1ESYK1lqyNzIzIrD0aiPEr75gjjjjiiN9THAnoI4444ojfOlT1l//X/9zc/MoCsZe+a2OIqkKESEjIyXfRhxSjSFJNhIxEAnd90/quH/hVVFUPmADVey9JDHH0wfe+7zwSWec6H8kVs0nRBWzamAbFygMrhrxUs5bLqphOp4CwXC6Xq+VqvRlYXcLMn6oOTDcAQN/lhYw1JlcUzEUFR0pCs79zjNEYySR13pGZAbRtW0OMiCqSLS+C9+nLLTj+Qe2ZaXFFBMjCYgFEAs3OEwoiWdFzYERBRKCgSQbGF4EBlQCQdGdbAZobWve5qVn/syM7Rm4PcZCaIuQy6/gFwEAmDtX/9nYeOlCQD80uHoqqxy9DOvGwxU6wrcpZ2fVgBb6zrh7bCXbVEQ9OdsiE7gnLXZfBfvG+o6sBAESESFVpcITIpOYBj72X18IB6Tz0wYEMemBVVQGscVBMiZImUaCQUhBNisi2KOt+vVIRkGQMzi4vse+btl3dXt3fvC4m08lkxs5FQBGdzM4uHz/bLG9jv13f9pPJ3E1mtnTGzFC726vXslWFpNPTano6PTlZXr/ZrG6Z4ekH346SQGWzWr599ZkzXNe1TicxStf1TX/97Nn7JycX3qfVsk1hc3f9Vk5OJpOpM7bxt12zZbZ8cmaq6cnpxWa9au/vK7/5r75x+au365t128Z9g+9Y4XcGSW59GUs44t6O5aB1x14cta27X+605ztTj4OAxcFRRun8Xu8/bv4lA+NghODYc8qIF8/OP3z/8tllXbhgLU7mlUBq220MbUipnp0r19vGv/zFLzDFs9NH9WTa9e3dzetms+TqpJxdltU8+HW3ul3d3caoZxdPnzz/5ubmum0aCb4sq8ff/E55enl3dfX25YuU+vnZh916efPqxf3NG0nhvW9/2xBfvXn7+uVLSfiH/+xPJ7OzbdNt+g7QzE4uq/ksxe72019wai7PFiJzMhNF64qyYPUdGAtVNa1ns/6+67ZNSMq22K7b7WbbtT2ofjFj/+uGd4jZfGtQVDUAE2vnZVlZLhgtgSEwhIYJVTSGhCn2iYTZgEQJrNYykTHGpCQhhKKwSMBAzMRM1pI1OftFARSRisIxMzHZ0WpDVDGBJLLOOWdVh1ghjUnzTMaWpgZAZkRiNYZLL7Dx+LNPr/7N//mDH/3y1V3rIw4M5pexz0d8ZfhHMLs76ev+FVBVCKBLnz6+TcVPX3gBZPP+o8WiKr33gimh9jHdN82r6/Xf/OTzv//47eerdh1SDyD7Z9aXnO3B5R1Hxw75SUNMhCLiQwgh9L1v23aI3hMlSQpAnMNvmpIY5hRTjLkgZMqpb8ZwTr1ipuyzAQgKGmPKeQ+DvRNBNmTLczxmzsw1JlRNyiREgyfVw9GROWhAsISlNbUFh8EAWsOMZBAMIiswkkEyhpiRGIEEUBEwJeh9SkkBICUxhvOsLz/6zKpRgBRTWRW2rNR1nama1oNJaOj/j4454ogjjvh9xJGAPuKII4747ePf/tsP/8V/88P/7X+Ire+9bJtV77sYU1UVRVEQmz40XR9DGAhoawwCxJg2q03btNY6V1jnDJIgCqCGmFQ0EYlojOJDJGuZDFjmcuImp0Fumi7KIKw8IB914AytNVXlyrKIMd7e3t7d3q02G2PdkIk5Gi8Myk3VGGMSAYW6rpyxIQTvfUqpLMushdlx0HhQclBEi6IAgL7vrTGEmGI0xiBR0zRZHP0bIBchzBqbgdsVBFJVQiQVVUIFYDbZqiLvNRLl2cMQEFEQmUhER5PlUbVLREhMSMS5gs4oVR4OxcwIOOias5f0QPRl6n5w48jXmgWIOzoadmYMeOixsV9W4+DPsGcID6XPuyACDlTmjnfMp9Vsy0iIuqsn+JBc3hltDPnROKRHj+WFdJTswsH1qA4UqQyH3Mmld2UMYfRyOHATzpCDpsuXJCGklACZq7q5iTH1TGjrgo0FQGOMq2qt6j4mV5SgqV3dO1uF1ktKeekbQ397f13NTpwrTVH5tj09e4KAt1evNqt70ETWWmeNda6symrSbrakVLi667qynvX1tt8ufd/d391UZaknp4S4Wa8+/fijs7PzyWw+nU5ikm7btE3LvBFFVzof2PuubbeuKKuq8mWVQi8i0ffee1sWCphSrC0/n1R/9N7F1SZ8/OY+Zb3eyOPSUD+Q9sT04Lwph7nJ+GBpPkQI8iHGyAjuO/cg2rDbZz+eYR8PeIeAhoOt4ddBQQGYaD6tPnz/6aN5xeKjpJPFBBl853vfhRj6Pp4+msQgq5v7ru0uL8/qqkqxv725ev36ZVVNz87Op/OFSOo3q9XN275t68ns4vSsW6232+3tas3OPHv2vFqc9pvt6vomxfj08ePUbpe3V22zLgu3WFxOJpPbu/urq+s+pG9/+N2ynm227XLdKPJ0Nqsn065p7q5erm7eXJ5Pq7LuY/JCgkzGtO3S960xjMb6JCGJiDBAPZmRdQJbUUAi/ULbfJ0xBKZAlREKoIl1M+csAoMSAAMyAEHOpFdJlFASJCajCpISWGZiZ51oSilB/pnJGssGR5/oIfEj20CPDh2gKpJAVTUlFSEAQkqSVBSAVCWJBB+MYWuYjZEgMaWoGJW98Cef3/zdjz/7dPsNYQAAIABJREFU87/5+U3nOwAZYyH4O9VBXy/8o1v+SzloAWwS+KQ/+vTKh1AVlvBbxbNzrxJBAsjd1n/y+u7vf/Hy+z9/+/GbdQMQAP4B8eqHHPQRMEYrkXKSlYjEEEKM3vdt2wEAERFzCF5UmE02EMva4WhCnqR1XZ/d2AYCWpWZEUBUiUgxs73GGFZRHLO9QCEEDzm/i4YZ1BBDJwJN7wQJcpaZDM8ysYwFo1EoEQtma9gZcswGmYAoz3gIgPJxNefqiEIUEJWQkkUkhfwWkFA6L6JJtAzReaUCvcMuxqpiEP2SpjviiCOOOOK3gCMBfcQRRxzx28flJfyrfxW+G+/vlo103nfed71vz87P2BoCaJp2udp4H1QVCUpnDZtMGxjDzGSMscb2fisSkKAoKuucYWPYsMl8gGNbClssalPP4aefbrZNTCIK8mWiPmYmMm3bBoHtdtv1bQgekJAJBSVzAyq5/Dgi+hBUFAmjDyCaxc7e+1zThpkzfQmAudpa9tlQ1aYZKOm2bVMIg2sH83+CAjqzEKKAIAKUV7gIIokIkEBVhAhUkihozhLN15BlxzAqoEeHZ9yrj/dpqKMWfK9lBhgtEYb80yTMREyDSnSQTeOe8hsIQdlR1QAAuvP93ZHCO4XsuFZ/QOEe6J5hV3FuqA40brajGnEnch1EibJfWj3QWe9luQfUsOiu9tABVz78eleVEg70zXuV9hfV3IenOPiDiCipbdvgfW4iIibr0BVkrDG2D+pDAEA2VolCiH3bkmC7WkrsitIaWwJxH2PwvSHOEs6QbDk9mYa+79um2Rb11hWWjDW2ns7O/bZPfR+aLWBRmGI2PTFEfd/d3F7Vk5lz5Wx+FoM2683y9s5YV88W1aTyPm3WG0BbT6ZlVaZQ9S10ncfVaj6blZOpoPZdFyU07bpmQraurMHGwrk/eH758dvVi9fX2z4d+KnAkPW8G80jhp8OOmtvv3HoqfHgk4yj5D8v3ndRiwN5KO5tUHbjacdT68EmD2ibnXX1eLi6Ks9P5//sO+8/OZkUhEgGTSFRNCaNqsBn52dVUfU+geLJxZPZYupKu21W3XapiJOTk8liQkbb7apd3zfrlbHlfL4oJ/Xd21fbbotFVZ+d16cXyfdXL1/1bbs4PZ2dnGzv3qxu3oTgF+fnZ88/aFd3b968Xm+a+fzk/Ol73of1ehOEpqcns/m8a1a3b19vl3d1NZlMThRiF1tFNM7ausLUAGhSYefQcFTxKVquFucXTByBytm94NfaDFT3XfpgsAghWKSaTG3YEYr3kdQaEkBBUqaicKUzzqAhsIbqunSFtc6wIVcWdV2rChFYa5wz1hqbiWYCw/lGCkSMCMFHhYQIKaUsV87jLYS4og0zO+cQMIn0fe99H7w3TDz4OEmMmsg1Qred/h9/9ZO/+/nLlQ8eQBCRCLJfzBeS94/4p4wHJj+AiASIChpU1l4/vdr8+d/+hxB823/jYlEVroxJf/X20+/97OVf//jz661vAPohVprnMUjDU1zf1UP/enX07zlEkgqpZtscy4NZmeTgNSqBiEpKMCSFqUhIKfU+N/JgrAEIADkIraKIIKLIpKApJhVJiccCt9D3vaqmmA7yfQBUk+QPedIv/RSrAkAUab2PlVW0jIZQ8+NIRAMkQGBQwJzhhjh8h2zIWLbOGEPGMBs2hpkYc/wXAYiHMLkqsMWiSra+Wa4CYDTpf/xv/+v/7n/6N19VhxxxxBFH/P7iSEAfccQRR/z2cXUF//Jf4v/63wuJTwmYTVGAIbJOFFMSAWRbOLJIaAwjAhNZ44pqCgrMxpWFLZ3vt6oBCB0bm4lPVCIgk1d0AVQ0QGygWd1t1ysRye4Pu5n+qMIEZuOsJSKJMRt6ZBIrhpCdJbLlHxMLMxGlmLLrRQ+Y7Z7zV1XNPHJmLJl5fFF2PGsmf2MIKUZJSUQwxt77+OW+e19clrwjaBrSRgc6bpQb47AYgb2HCIJmIV4m6mhkZx8caM8wj19GThpgoAez2vrAzlKHVZaKKiTZkboKgqN4ee+PAKoqiKgjCznW+RtSUA8vSUdP4Py+d0URHzpdICCo5MOO70T3dRn3Zwc4XOZl5fWhw4MCHJKRIxcqO3cRgB1bDjuJ9EO2ck9AH17rF1Rv+xMhAmiSlGIMse8AwBjL1gIbZkNsIQYBQCRbFNQaIEZiBUmxj75ha00xQcP9tgeV4Ls++LqsBMlUk6le9F1ze/W6b7eGWcva2bqqYDqdh7YJXQe47Y0rXTmZnAgsb+/eKsBs5opyMp9r6rumWbXN1hRlWVWhl6bzfd+6wlZlwbDYkmm7tmkbZq6rsmZUwu1m3a/uFA0Ql5MppNDF9Oyk/Naj+Ucvq/tX92nP2OfBM8rK9yNk304HDXvQeIdN/sVcc9UHG7z7IXqHW8Z3zrfvsJ1KHh/sSYyzSflHHz7/g/cuL6e2clpUTtFKSAa4sCUAXzx+GrxE3xtjJ9PHVUUqbWhXkvpqvpifnxvHPmyb7XK9uovBny7OJ9NplLTcrtDw/PRyfvlUTbF6+2Z9f1NNZydnZyHEu+u37XZdTaazxakp65uPf7m8X9qifPTsfTR2e3cbYywni8l8EZO/evNic3vtjDk5eVRUs7ZbhZgioLHWWMdlYZzRVskwWYuExOyqqpotUkqujraavGuW//XB+GHFnUYYx/ASAhCARaytKZkLIgtsGYwha9Basoay2T0REiPlBPmkKWqIMSVQgfwPCZmJc2YIE3MmBXMkDFXVe5/T/VNKKkpjsUsRzeVqjeGUJMYIoCKSJBkiBBTQGCUKJi5fr/qfv7774UcvP7tetgAJUAAJUPHgNvKbNtJDfE17++sNHUPAQeW+jb98s3bV5xHwT7/7LaZwe7f825+++vEn1y+XnVeNgGPVQdzt/ZB1PsRR/vwQ+emxs2hSVVVittYWZbmbABmm/NAfqltrdnpPh9Oew+Q2IlQFRCFERVTKsXOVlHLfptHlOZ+XiA5mVKoqX/rJU0AFjSLbEO6bDlKoUCrCktE5Y5kcEzJnPXe2+kGGfOMy1ljLzjIRGCbLzIhEwIxD4J6EmZmtSgJCtQiTIkp924UttyYeKZEjjjjiiK8Cx7vtEUccccRvH//iX/zqz/+XsizqqpIeDCNlaTGhKsSYTFHPyhkSG8PWcd/1oFBVlTHOsEUiLhyXFlIHmoBRew/BY0ohdjF1g/uyDz5IUgNUbm7edM1aJCmC4kMFEgAAGObCubIsfWpzaZpccC/4kESIGbLpgsigHR5XDjHGBENWY34PIhJjzJsRUXadFslV0QfjixgT5Np9qkgkqiGEGL9UAf2ljMBDBo2Isu/HQLdSdsLIWzEPJQSBEAhlPKgiEFKuij4eFAmRx4TxkeVFpiGBfPCdEB2lxTt59CHNu2exdac1fSBh1tH0YzjtTqelIKO4eTzc3vzkgBbfN4DmIxGhiqjoaPA6nHtHOQHsVn+DOwcMB9bxaumQFj7w58heHAI0HnD03EBEUcVdRfuRid6xmQdi8h0BvqdO90w4IYgCoiTpuxZAkQBUNURFVMCyrCbTGThHxM4VRV3XdSUxWcPLvlPfZ+YsxDA1M4n+7uYaz87tZKpqrNSL08u7m+u+7VBUoxQnJTOdnZ1vV7xZb+N2BQA4Py2rekLzm9u3vvedaaZTe3p2ShDpnrbtNt7dXl4+mUwmxhZt263v7ydPn1bzE0JWwK5vV6uVtca5whVxtVptm4Z4VdYTay0YultfOXAfXNTffnr66dv7NooCDi09dvVDx5J9++/DGQ8+ALuwxcGrO9vnBzv8Ok5t13GHh90f6sFu4x0j85eVc+89Ov3nf/Lhec016aQqJ4tZ9L3G6NiaiXWqpiiX929821nj2DAStKv7frtiw9PpeTlbSIx9u+2b7XbbWFPMpnNme3t/08V0fnZ2+uhJWc+26/XNzXVZ2rOzhbH8+tNPr29unLWnp/8ve2+2JMmRXQneTdXMfI2IjNxQKFQVis3iPmRLS8+IzIfM7/Q8zb+wn+apX+dlRFp6ZHqkRbqq2STBWlBAIjNj89XMVPXeOw/mHuERGYkC0QQIsPxILu7mZmqL2qbnnnvuk+lovH779vrqSiS8fPmDFy8/uLq4btu+qseT+YzQf/mrT66++O24CtPZuVQjJzGHVEpxR2bNiQBEokhljuAoEppRM55OnKhdd11fVG8FfN8z7GI/uLte70ijXZYEsENkGsdQMweiWmIlWA0EtGAQBPBSCjkRkIL3vZZSkCRrQYQqyu7e4O6uZuZmLBSC3CVGuA+aRxIeMmAQgIDcdVAwhxhFgqnmnHIuo3ETY6A9NWUAxaE4JdJfvbr+T//1k89XuQUY5M+OqDtLKAAAfN85/hWO0zs4ctDfKnxnS4WE7O6d+kULv/j0si3WzJ6mvvvkl7/++SdvX91sNztGEgEYYHiUGNx6Pb3bm8eefBQ7xt4BYKgULcxVVY3KUIcPVRUHH/cDv5TBUg3uP2QQcXBaAwAzV1USRoRCzEQArqUgIDGXnAGAhbWouyPtPMGIyOx9Nvs4XNnJbJ0Lbdq+wxHaWGgcQqNYR1Ih2LlXIQ9vrYyEwAzCLEQMCKaeVTUDgiM4AQypcaAcQ2xGiApICkDhbDyKV31fd3XBr1mS5IgjjjjiiH8UjgT0EUccccQ3DkT85D/8H3UdT86fMMzRFIkgBnQDMwd0isARihI4Eoy0gCntGCsD8NSudZ3Re3B1N83F1YTRsThk82KlaC6bTaceq1E1lHmyLx2ns/B8OpNQn55cF7W274mlqDqCiLi5mZr54LCRczZTAGAiN+/7nogGk2VVzTkP6rZbBXQIYSCmByailMJECOhmSDSoY0rOqf86x9PNdE/XDoYOd54DCABgu/pWB4YVw5Lk4Db0yK4I1jDoosGkEMzMTIF4YKVpV28L9rzqnqYelNa7QoKOew76zrMAYE817k1YEeBOeYp7PRIB4k7UPMx7y40f8JK7te2oawSAoczO3Q77Ha14v8cf2C/gncDa7XCdvs9p3kkmCff7sD/mex761gvksLbd/fU9wgv4/rdbVtzdzA3AwI0omPq6X/frtSPUTVPXFagODpJEpKrbzUpTh4gcQlVFEFqs1g5WNVVVh/VmJUWb0ShWNU5mH3zww5uLL9Y3i9KlOob5dFaopn5UVpv1zRthwNkkROEgdT3fbJa5v0TX6vx8fDprtd+mvl1vrvHyyfOXSNR1bd+1y5ubZjxRAIkxurebdbttYwhNMzk9g+ksbdar0rWBkEXA3fP6bAQfv5z990/Hv3q7zrY3wvZbtepBl991mz9QM9/n8m+P6C0X987hxvcM7++m+71WfxcI4Ml88ocfPf/J81lDSUiaipsY1u02tRnY68loMqo3m816ubCUqumsruj64lVql+o0np2cvPyIqNK0pJyxqMTm2bMXo/G071O3TRKnp6cvR814s1m/+ey3q+Xipx//ZDqKi+u3F29e94U+/NFPnj47z337xae/EeIXP/749Oxpu22vbhbjyen06QtmevPpJ5/84r88OXtyevpsPD9TrpQkNuNx6rOBBLxZXFHuUl8AGBQGK9HSa9v1utP2g+udC/f3C7dBpIM4wk77DO5gMKqreV1Pm6YiQbeStVfwApmRCZiN0QkM3QKBMITARIzITkCEQtQ0VQhi7mYG4CHEncQQTYRijDsJNZOIMHMpRYu6WlUFCewOLDLUpB1OcjVloipEYgKApMb1KGP4xS8//2LRvl3lTbE8sM/7m+jRfOP7iXdvUcOJae7ggAp+3Zm/Xtn/+3NL5ep6dbXtCwIObz+A/hVDDvgVb2m/V/Adc2/e972qMXPTNDHGzWazM9TCBzF4QEQSDrJjCW456AMFNAGA2s4WRU2HWhghRNgnQ9jg2hV26RG3b0e5Ry0Kpg9iob5/Mjm4mgIJMROQm/V9KjlvARhBwAJDDDSqq7qKIXAQFiFhrqLUVawiB0YwlyjM6K7MLFF2XnZBgtRA1CMbYjbLeTAfOdYhPOKII474NnAkoI844ogjvnH4X//1a39VOI+bihw9OYC5ZzB1UzVQyAY9Opg7oCOYW0mlmJq5A1BOfepahAKubprzQPIKsBmqWnF1UNu02RBVtMuay+Ck8PiQjJiFd3nXgxzGEQFJAJBQRMzM1MyMeBC0saoBgBDBUIUPcSh0bmY5570AeieiqapqIKaHoaaqCjHtJTa5lNVyufNE/hrHEwD3JsUHEw0Ga0k3cDCguyHrfuxDAAQEsDNbxjvaZmeKsGvddxYUu4VhN/7dL7H/sF924G5x//mQyd0zyoPu+FaK7gfGC7cc8V4V7Xf88y3He0d/734xvKUwd0vdc2jAB4f2kNLc7cOtYvpOBT2UsQPc792ehN7/4jsjyJ1/h++36H3ddK+ZXbODDbSVUgwQYlVvEbIWtgJmbdeCY2iAAKzr2u3WVGsijDEVzX1uRuNQRTNbL9fmCmboFgITSzF1K+qQUprNTyx3K3cteX1zVQlzaKSqq9F4u1m23QavL3OxWI/Ozs/drJSubdfXVz5/8vTJ02cIeHN5td12crOYzOaj0Tj1+fLy8nmQWFVEEcHAmxhls1mLxMl03m43V2/fqFBdVyKj2WTO26Wj/asXJ1d/9gc3//HnV5tUbsMLj1yWDxhhPzglvhJZ/I/kXr7qvAgwHtV/8KOXf/mzHz+bhDrQqKmEKHdby8m0UKxCrIilX6/6lKZNPZs01q2/+O1vJFAzm8Z6GqTerFZpeZMWC03p7PTJZH66XK8Wi5us9uz5y2oy1ZTbxU3fbs7Pn9TjZrtZXbx+1bfbDz/6ycnTF8v18otP/2G9Wr744AfT2bzr03rTPXnydDSeEdjy+vLm6u3LF88/+ODDuh6pAwJkNQEioJzS6mbJEupmDCW3297dc8k5F1NDcC+5DqJCiP61tbX/vNi76cBBAgbAnf4PapFRCBUxuOakamYELqiGwiAOTs4IBKAO5FDMBYERhYf7thGxSHB3REHCEMKQNIOITBRCoOE7ETMjUSnF1MAsRGHhvcEHESILMVNKCQCqEIjIEVkhc1y3+svXi19fLBdJOwA94NEPdvaI7zV2ITZzv33QtcXLOvW/eW3qKWnZUc+7+RHs3SqpeO+pecR7MLzpOIDDUA9iuELdIeeMNBQnBLDdI/2WgSZE3nOyw81lsI0a8iD2hmeARACOBoPrmYgMqwAAMytahuUdfOfYDKalvNub+xW5g5u7aSGsqiAT5ugqVhAc3NAN0B1czVPJQK7GqRAREkIQqWKoqxCFmCD2TASlpFCFqo6IyMwxBiZ0xIyctnzT5a5PKuGRPMEjjjjiiCO+ARwJ6COOOOKIbxw36e3z9cvfzD8pOcW88ra11Kn24KaqXde3XUnFQ6hIGHeiWM0lqbkDEkvOOfUtog3mfDmrubOIoRVXNQckJikagKCHvNjkTZvNDjS1B0CEEEREttvtZtt3XTcYYjgoEKLTkJU5eDQzDEmau7zLwbPitsbgnnOg29z1EMLATQw/3QqiGXeVpm5Z8QdJ/18diEjMe9Pnw5HMTmuD4Ig+GAUeLhiEhcNO7rhnXMHdgWA3QLorEXfrmmhme731g5X5u7JnONivfet+V10QbvXY7nvZ8X6f9n4XhztzqLy+RyHvlciwL0V4MIPfemzeMtGHYttD3A7xB88F31HvO7H27Tb6rl7RwV488HN4V8i7n3q4l7eTTVPfpZSGvkSkofFKYtclVwNzME8pMyE4uDoAAjMxhaoCIthuAwmaa86qpa7rvO37dkvgWrIIjWYn7rBZLrbrFSNNTs6Z43g6B/DlzfVycZVTP5mdzc6ezc/OVjeXfbcxtRBHs9nJbDJP27RebxbX1yJRQtVMZqvVYrG4Oj2ZB4kaxTyYlc16LbGOzbiqRiFELUmLxlDNZ6eMbrY+r+1Pf3D6355O+3Kz6orBPt5xjzS5J06+3zcPL5L7qufHhvEPO/kgDvOl8z22HifCD18++4ufffwnP/lgwl5JCLFGoLxpu/UaDCYnMyNfXV9tNuvQjEbzKQktX39euk01fjqanjWjOZSUVteryzd5u61jfXJ2bqbrzXLbb0aTyfz8DAFuLi4Wl28roSdPnnjR68vLzXJ5Mps9/fBD1XJ5ebFYrebT2enTZ6XYar3OBV7M5kRwdfXm9esvVpvtBy9eTsfjlFLWNG7G4J5T3m63m00fRun8fFaTJgCwIjIo9IA41FWtfZf7vu82aj2RP06NfLdxG6h6EHNEAAKPgDVRQAQtKaVcMgN6YCRBJiYiJgkUAzVBgiAzIliU0NRVDAHAU051XccqAPhQhNDNmFmChBAAoJRCRAhD8QAFV3dnoSBVzp3mEmPEgVwCYkQOXHF1t5lIJHJxs/2bTy/+89/8+pPXVy3AwEIOORu3kTd8/KQ/4vsCv3v47yudkiOAZ/PLtvi+tuDuD/qePkWAoUQewO7EHoLJB1T1kYd+BwiIzKAKCCy7tzIzT6nfbDYcwlDb8yA96zZPav8MOJguTOZu5jK4v7uHGACxlMGEg9x89wq1K8hxEF5HJETznY2ZvxMy3cfsB/cPCACTGM7HTQ0WQIcQPoAPBLK53b5LFVVNxcwAekIUxiAcA4OpltynVDVV01Rd3w/q75ySgWPdaHOTOEI9khHwUQF9xBFHHPGt4EhAH3HEEUd849h6udn8og128eYt9wvvWtCEPnhUlJQLSxVCbVr6vu1Tz4LExELD+/VQgjwEKZqJKMS6dkIiFgECYJBQAZA7UJgoNH2J297fXC4RlQnKY8KOIIGI3rx9s9x0i+Wyy6Wo+V5ulplt7wDIzKaact4VGzQjxEHafMsvq+ouQdpdRAZL6FLKbZlBd0cHGgQyiKnvc85f3291MKeGgYqmW+0f7LTRhkho5nqf50MoqRClwXzi1sgZwAkzEu3kN3sWeyhkCAA2FMy5G1Ld2R7fWnPsvhwooGFPtu5kxXC4MbiXG9/tE+4NXA9Vr7uPd74Wd5Kvvf7LDmj3W6HggYL7nrT6Trx9sLWwP3R+uyTcFovfOWHvlNF3LQ6z+cMown1p7y37/ECe6YSWUuq7VJISyuB3wsSTZty3fclF1RyAiEIQcrCsRBLqxjSre0ASYjBDRDPXUtxUCNW0aAErKUPVjAFJzdaX3fLmhrgez06aZlzVzabt8nbVby2IlOm8GY1y36WUcrLVzaIJdSAZj6el+Gq53Kw243lsJpPi2q0uW8FmPCWWUIV+2+eSUi4SmtPTs9n8dLW87lPKqVSxyrEJuK0hfTAOf/rR0+tNatMq7R0eHg697wvUvwR+79y4+/aexQ57+Hbmr8LTDFo5nE5Gf/aHH//lH3380bMT31yHGEOsCNxSTtvtaDKWiktJi6uLvujZ8+fVZNyurhbXF3WU2cmTyfxpCCGtb9L6utss0TxWs1hVV5cXKfexlsl8Uk1G64vL68uL3LZPnz+tY7i+uFhc3YDTy5cf1E3921/9w83NVaybFz/4kEN1cfl2tWons9NYj7bL11dvP1ssFvVoPj99ktNms1oAxyCcc+67brvZ9n1hksDBUqd9h1YI3NTMgCgEiZb7brPMqXPP71HmfS/w8FockiQi0Vi4Jo6IDCBBJDAjBeEoFISCIDEMtQeBkIRD4CgsjEwYKyEiCYPfKkrgEAZVNIO7mebsdwUMiUJgNTOzEHlI7DdgBAhBiAmJiGBIhpEw/E5uUAw7w3/4/M3/8/O//Xy1bh2AaH/bub1pHvEvCvvHJO5dfd3dbPB8vqWc310IAA5OBtyd59/PzIVvHg4Opg4OBrlPQzTdd7d3kiBEZKoGgI77mqW7x/StH5HfPrz3r3lq6u6mpu4AUHIiFhYenvluBkN4nvk2kH+7RSUn1/v+G7e/7cIT4OZIBIgllwKK6DvJAYGaOQHgrgYJIVZD4oVwYBFhJhQCZmBCQnAAZiKmXAohxRjd1NyNRZtxC3ydlZEfr4p4xBFHHHHEPzWOBPQRRxxxxDeOG9sWHlu6XK/XsF1A6smNmQeT5WI4kqpuJrmU4mCewYlIQlUBogGY2eBdl3PPRFVTMwoRkxCiE2FV14Ck6lJNs1U3G+iz3ay29tCmYgACuIgQ0c1isVxv15tNv2P8cMdRIu1GEYjMxCwpJTMDBGNFxJR2HtAAYGaqZfisWph5SMMcCOjbZMyBLhxcO0opOaevTUC7OwzL7rngPd/rsEsMtUFT+o4csADQXlp1J1/eV+iDPVuKCEBIg4D6UAGEB8MzuGOFD4jZA1Hx7Wz3xMHviIT3TRwQ0Ie2yodj7ftN7DlkhztmHPajyN0WD8dr/w8A+mHb7xLQw275btP3KdJ7Wdohx32v2UPco1j93vJ765LA4GZWtOt6UgdhIhJCqmpTs5RLLmBeV00QEg5DFaFY1X1rbdu33qU+azHgIIEIqd1uZ/MzAOrbdbveZrO6GdWjqRW1rltd37TrdQxVmEUKcX76pCXU1JXcbTfLZjRtxmMDXC0WqevXy0U9GjejkaozcJdz37aNyGQyJt1u+zaB15NZVTfkmrq0XK2vLt7MZ7Oz83Nzu7m5ubh4fXZ2XtSIuBZ0T3/5Bx98erW+XLd5m75kmPtYusKjsz2gZg5CCrsP73Tv+xZ9PxAhBvnRD178m7/42R//9AezMax6rJoY6xpLGa6NJ+fntchmvQZTRpyMpw623mxyyaPxeDp/Eupx3202N1d5uxHiZjyeTGbdctlu1iJhPJ+enp07wtXlRUr9dDo9PT3pNqvLN29S189PTp88e765uHjzm18nzR9+9NHJ02eff/rZm9dviKvzZkRV3Cxv2tV1E+OHP/zo5PTs81++3qwX9XhuAOaecu9aqhgnk4mW0i6uu+0a3VPXG2pKigyluKDHENxNhL92WsZ3A74vRLj7SgCRaRJjwxQQGT0KRyJhEuYoJAxs2IYyAAAgAElEQVRMQOghcBAiBmKSILEKgkBgzChCMVbuToQhSBBmIYRdObLB8ohZiHBnAG2mqsw0hAMDChEEYd5xSI4EREBDZTBEBWz78vnlzd/++vO/+fWr69bTl0v8H6cmv9rxOfLY3yncPQMREH1f/PQ2nnx3T0Tf6eDvHrxHyvArYDAlA3RwLSWnlEsGGIJGxMREOJSr2Gc/ASAO1POtrdjuzWdXNGNwEwMfCpLuChIaoIIiAKgWLcXNiEhiNRjsw9C+G6J7UfDH+N6DVyQzKOqpaOeOBEDgiMw4eAQ5IN9WHSFklhCkirGqYh0jEzA6ogUh2d12AMDVnZCEmQkBoQD4aNpSaN9eJYcffXZ5vDscccQRR3wLOBLQRxxxxBHfOJQBDEhEQkzMGBtAQglVEGIGx6pq6qoZI45L6fqemDhIqCIAAAIycRW5qrxkRMQgqDZIw7AkKBnJAVECAXFfPCUtxdUglYfy58HrAByYmUVUNeXcp36x2uRiRIO0DQdFMw2OFESIlFJvZkycJAFAznkoOGV71FWFiH3qBx0cM9uOhmB3N7NhoNO2myEDNOferHy14+fvjDTxVlXrtx4Te2rUFXeWqHfC4dulEMAOW0RAoN187nirVX4nPfRQPLrPUL0VGx/OcLvNOzL6QGh9n4iGgy+/U5iKd3MdNHVQYvBuRH4wbb+BDl82sjpYOe5p4j2BhbfVEB8Ozh6Knx9niu4cOgbsE6h5ZzzZt13lGmITY6Vdl7qOWChEqiocjbIqAQzp+aZq6CIsMbjpYrEo6qpaNzHGsFgsWCqRgEjNaPzFq8+Jw2QyG03npc99l9tuQwtDsmpyNhnPIadV323W6yqOlUOcnNQQNm2CvFmubrLraDKfnZ3knDGnvN0QaDMZx3q83HguzmoNk8TJaAym0HftxZtXT1+8HM9OUtHUbrbdUqrROJxRXeFy8TzIH/3o6Ztlt/r1G32sD74C9XwYR3kQORim3mrnHb7sXHr0l3uND1+DyPnZ/H/9t3/+F3/80ajG5fomNlXVjNw9p76YTWYn4eSk3WyWq5W7v3j2DFTbdt1u1sn82dlZnM+NQ1rl3PXdpovNdHLyPDTN209/lVXHZ2fT02cUm+Vnn/XrdYxxNJuCyPr15WZx3YznT17+0JrJ9S9/CVlPT87mJ08urxavXr+OVTw9fTodjW27TdsNmZEQOKJIVcVFSV27ZRFVK7kguBCs19elrnPukqaiXhEDctNMqjpMJ/PUtYhEJAD8Pa1BaLtrHYgYEF0L+s79OTJP6qomCmCEwEjCyOxRoA7EDEQGbk1TV1EGf5KBGiYGQQIohFjX1XADIKIYJARWNScUpqGcKxPBzkfIg3AUTjm7GzNHIaLBT9bBTF0JBgrbTL1YSRbfXK3+7//0//3i1xfXW08OOtw7BtOFg/3cE2IDBf01yKJ3HyXfWXwVQ4Dv0e7c4qDj9s9DdUdXAPR74d3d7t1lN91lEh0w1A/vh7/neOe6QL+LQ7tv23a1XgECCxGju5kRwD6ADT6wzEmTOxDTEF6i3ZsgDS9cPATmkZjJCRExxjCsV92QAjFrUUIMwkV33tNDthwMbDcSgN7rtsNHmqM6rtu+AgxNBTGgCIqQIDAADncn3NWKBjfTlMxNyS0iABigMasZlgIFPIiEIESIgOxYS5QgToFnTQ6TV4t1yf3/9n/+x2+4a4444ogjjgA4EtBHHHHEEd8CTIM06zAez5+c+QiAhJAJiSUgMwCJgzgisSCE3fs5sgi4DcmM7mh9MVVzszYNomK1AppAk+Zkrg6eiqw6ulzTYrFJGR5VGO9Eu4jCGGOYzaYFWB27PjFLDFGE3aGUoqpVjIioZsI02GsMSpkgHEIIEvqUSiluVlUV4pA0SSIcQlTVnNNeAe0IjgjMDRHlUtbr9T+N3OSOBfU7FvZ2eHpLX+w4WHxApTo4KADiA+GjvyuWO+BpD1jVQ7nxfWrZD3/YG2a8bycOCMT309HvENCAdwvfrv9wC+8avfNf2B2KhzLo28Xu6Qt3e+H79u+Ja+8ds8fUQw8O0N12mQMgsISqipx7Vcu5lJSWi2Xb9aN6TMiIFEMcvBIYoYqV5g4AmZlDmM/ni+UGAKwUU23qxt1LLjFwrJuUctf1EvooYTI7uXzzmplz6hfXVxOXyWQ2nszcrGs3piX3XaiLSGhGI+1K6jbr7QpEzk6byXRqZiUl0JK6lkIMVZNS323bUT2q6ylTAAezvFkvJ5t5PR6fnZ0tl6CuVjJLnEwmleD6zeWPn04+f3ny+vLmYv1lIujH4O98feTC8Xc+fK32d5+J8PRk+pd//rP/+a/++HxWEWRpqqdPzohku9q0qzW5nZ2c6rZd39ykrq9jVcVYNFtO6qASm7OnEmjbblK7JkDiOBrP62YMACQBilX1OEjdrdZvXn3B4PMnT5rxeHF19faL15OmOXvxPDbN208/67bt6enp7PycOFxdvhaR2XQ6m02R8LPfflpSNx7VcTxvRiMtGdwAgJhDqNyHoljMMahqKSnGkEVS6seTSTLIphIYAd1Ni6ZUSrZHlXnfG+C9yw0BAmHN3IgEAAYgd3RDp0AcBIWBBQmJEIRJmFgCM7Hs0kSIXISY0YeKtjiwWObOiIOnK5qru5k5EblD3/UhhBDjkIZCCIPEMqVuKFkIbo5u2dWzE2NoVuv+84vlP3x+83bRJQNFMIBHrbgfjfUd8S8Ad08tP3hMPRZpe+/3Ix7F8BDex8GHchTTyWQ1HoUQhpCt3VV0cCLcmWvtawneZYftXgd4aHhQRevulrtTNoChuzMRI+EurIdGZu6ECMCAYFqKu6u9m25ye2GbozplhW2XNeWWIAQSBmEMTFEoBo6BhYkABmtrMO8RhSgworjsNhIQkYUk8LACBCQCIjQCZvEYgpBkAYCf/8mfwC9+8Q32xRFHHHHEEUcC+ogjjjjiWwBXpbt+OTtfz0+nGDLGCpDczIEd0Q2gT94nM3URDgHMwE1L9pKtFLWipZSi5mZmORciAnctGVHBc2q3qtlN1x0sOr5s481ik/MwRHh8mEYEzBSrwFWNUvdZt20nzHVVxxBYuN22fUrj0QgAcs65ZAAIEtTU1Mysrusqxm3bDm7OsYoAWPVhMBaMsSol912PRINThGohplHTAEDXdddX1/hPWfXFH1eR3uPWfCeeeWQs+/hRekysfPDlITH4LlE4AB/RJT22rlth2GOtHzR29/GewNgPSe5bqmbv0wHvCKEPPvojn+DhHt2OZG91Zw8WOiDFH50Bb/fS3Ya2iZmNEVDVipkjmTsQMzMUVfUgAYkQUGL0kh3NHcwckcaTcRRxNTePIeSsEjhIZN6RZcNKiSRWo8h1SW3bdXZ92VSVhNBMT0jiZnGjtnYKXI+Eieumz30uqW3XaTyZncwcfLNapZy072KIQYLmXFLOKTc1VfVIS95ul5vtdnF9QWihrurxeLlapc16MppMJuPIUNPVB7P4Rz84/eJqff23n+vvUCj/Tn7tG+deqhh+8OLZv/2rP/3Ri5OKNBCMmnFV1Tml7Wbdtu14NGpm8/XycrteA8JsPjfVrus051A14/A8zE61b/vFVb++RrXJyZnEqu+Su0nVzJpxM56YlvXNdde1z87PJ6NRSunyzduuz+dPX8yms7Zdf/HprwLB2fmTejwp7iFWdV0JD+XuaLvdxl3wxZl5sJBt6jqMRqqKxEQ8kKQSQlWPMJUQY4MsQfq+AAExAXrJCdEBIBfLxd53N/gO4y4LZJd34YAAhFgxV0yRSNwIfPcHXRgH5w1CYMIhPYUAYhDiW+chdwdmRIJSMgAgIRK4s5k5OBMys+XibkaEDu7W9525Ig1e/AhoAOSmKfVRhENAdy8lWy5QQCIHentz/ZsvLl/dpGVvBcDwS/18h3yV710XHfGPwPscNt7znDrid2D/TEFERGGpmnrUjIKIiCCSDrwz4GDWAQAYAXyQPSMAupoNrvlw28wAylrcnYhgsEO7fQXZ0dRABOaupiRIiIBQMlrRwbvjXQwNmMNw905ZzXLvGdGJXQjqEKogVeQYdrLmKsYqBCUcqiVXgatAbiCC7MSE7GiAtiukDFld0RTUshXUrA4A//u/+3d/8vOfHwnoI4444ohvGkcC+ogjjjjiG4c5zH/4yrqwff02r15VdQWIKaecNaWS+p7USD31yRxIRJgdIOe+7dqcEzMjECJVdU1IqlaKAkCMgQWI3bQgOBHVddUalmUuZobIQkUd1GFfsw6GyjAIIUqsgpa86baLTQqBJzQCBxEiAgIIwgghCLu7G4lUzBxDzDmXnB2gijHE6G4xCgJKEHBITCwyeEALYWAeLDi0FMCahWKsckqdOX59H8+vhTuB6PuGrgfT37dl7yek3zPRD1nXA34YH7K1dwsfTr833t4bVR9OfLihD1vw97HidzKzW6Xhzvh5tyzeX+CQTN/P7fDoQfBD5+mDRfai650W291VLasxDM4wCEDj8aRtO2IhYstls+3OTuciwQERmZgHJWbKqW3b0XjKImAFdjESjLEREdXOHWR/HuaUp7MTQmu3pG1arW4m41GczKVunPji7dtUSgGvNVX1COtaUq2uJffr1c3k5awZj1LJ2RTctJTAbCx9LqVPqe+a0TjUTWzGse+26wWhTk9PQ9X4puu3y4aZphPj0MTasXz8bHrxkxf/7ddv1kn1vefhV7ws3uva8q7SHh/pv9vOetgWAiDifDr5+Ecf/E8/+3gSgDSFWNUhpq7rtm1OiUXq0RQkdn0yLU0zGk8nq5ubdr1yxGY8rWYz59BevWmvvshtRzJ+8uxFv+lWq2UuuQrh2YsXXIfV8nqzWlRVNTs5BbXVxcXiejGZnU1Pn4DZ5vLtenX99NnzajQGYlObz2Y3/San1KcUG2kmU1uuUkomvekuobuqqhCrrmslREQ0MzCv6qYZjdu0JOFx1QBBMTU3B3NwLTkKEzEAmdr3WF7rAODojgAEIIhNDJHZSnF3JOBAMYY6CiG4WQEDRxRkYtVSCoggADq6gyEBOuRC7mpmzBwoxBiYGdCtFHcCHHxdMcZgqqqGhKWUtt0wD3bQSAjDDHUVY5CSNOWU+0J1LC6rVfvzT37zX/7uN4uUMsCXxmaO+H3G1zNd+X0HIiLJ4FszVA8spUjO4M7EWtS9OKLvCGg3s13oCBCK8q7O3/AvDppo3xcWNDPaO7Uh4lCW0P1h5h0NWX04RAPdjVnENN+bEQEcfZASODi4MNVVmFKMWAkoYjEvbhpZmMkNU8opuZuKhBhCCLyLNw4xNjSJHIRFuK5jVVeOIMwhhqYOSNyrxy6U2LZdSeAA8Is//VP49//+W+uaI4444ojfTxwJ6COOOOKIbx7SLW7gpMntet0uFqkVJFTTlHLf9Zv1JgBGlpIGmoCgrogJVVF7tBxjzQgAwJYRiYlCIEAUQQ7MgZAqMzNz5vG6aJ+2Wc0AdrZ+96jVoZAcBgkhxJTzdrtdLtckNQBoKaZSiBCwaBmGIu5eVAdbZy06WHMAQNFCfTf4+iFiUXX31PcSguhQIV3VNEgYaCBEAAUtJaXU9/1QpuZbOv6/m9Lwh98e0WC9z0PjEQeD90/5ik4J786Ge674kEv8kkYeio7vkYyPp7e/h2t+B+/V1b93qQd+Hz6UgnTwVDJoilUIGBCZQ+WABuhI6tC2nc1ngOQAZoOgcpB9oxve3Czr+bypgxPeXN1MpmfEVMxyysXMHd0gl9R129F43HVdNjaknPPF5dsTCrNqFKsGQwNQcumqIqN6pixN0xCopq7drq+vLlmqWNWIBIib9VqEsYpaStf1LOtYhVhX07NzIFpevmo3axQ5nZyMR5Nuscwpt9uOq6ZqRqncPBnxv/rg9McvTv7+1fU26bdGtP3OFT04g6sgH744/5OPP/zw6bwqCygJjMC078vb16+bZvTkybPJ9KRdrbsuxboZj0eWc7vZllIohNiMTs6fbi9fry/fps2CKVSjcTw9I7pZ3VzcXF1VzeTJT2tL6255qaWbTE95NF68fXNxcaFFf/yTn4rwzdXFerWYTUdPnz0lYTMjwJJ6dMsp5ZRJ5OmzF7+5/I0BxioCWsrZAbs+Jd9UJ1Zyn3NfVCNh01S5pKwlqzpaXY96pW3b5lxKKSzUp85dqljFEL9HPNddmOj2luW7OrIEwAi1SMVMDgROgAwoiELE7Ag7WyQatOIDhwQA7gg+JOIT7sgmJgohhBBoqHE4sFSwN+/AwTmWkZB4MIrFGOPASbkbAsQoROCmg/U/S+DYLLb933766u9++/bTy9WmQD6yz0cc8U+KIfkJ7ioDOLhr0Zxy6nt3ACQiNKfhPU1VzUxEAFzVVPflmgH2L5TutxUuhtcGROIhhOyqigBDGUNEGGyjbfgLDgoIrlrM3rU6uk0U27HQxBRjqIVqtIBGFADU3ZiYcefm4+5uGiTEGEIQBHczBGACZmRGJyzgvYLl4Y1YMeVtRwCYHKPVGktfMjLDEUccccQR3wqOBPQRRxxxxDeOlJHRW03YWdd2XY9CxMKqWor2fY8S6hDrpgYAcx+Nm7qqiDmV7O7j8ZiQtFi73bp7iHWMEYlKKSjMMUjklFK7bTHOYtd2KSVVBSDc1zEHgD3tiICIICGGUHVdattuuVyFqjhg6roQIxMPgxB3RyQAMzNmAQTTO8p4mGfHWjgSs5mlvh+GAjAUQ9dSVVFEhnKFhBRD6Ltuu92mlNQez8H8TuARI4SvInn+nY0+OuVQbvzALRoP//O7rnxoWg37zt1PvmWTd+wzPtgf3JdIPJRND00/ost+eCzuGXE8aPgBM74/kvcF0w6ELBKriD2paYV1NZlCvzEgIGIJ4DB4cyMi7DP6s2pkqpomjdNvP3+V+j5GzikDumoBdyYyZiJk4hCDEul6vdpuxqPxi8mHm8nk15/89zbluN2Gpqua8csf/nCzumlXV1232qylak5c1dVKKjm1qdXZ9KyezDmOF4vr1G9K3sZmND6ZdX3P0YpupYnTp8+3xUK3af26TX293c4m0/Dig75tu1TQ+snJqYJZn1+cyv/y5z+62WxeXbfpf+j0f++J9xUjG+8DIT49m//rP/vZv/mzPxxR2barSRNGdRTU5eompX4+P41BtNt27aYvNptOQ1WtV8vr60sZT8/OzmbTSbm+WH7xmfU9AYdqfP7iZbe8Wb79fL26iIIfffRhyHl1c73dLAB1ejrPfSqqo9ns5Ml5CHG7XS9Wi6z5/MkZlFLUikNxA1PQwgCmZbvtAECRKAQSQcS6rq7N2z5VXMcgbdv2fXKAIFI0xxiIoJScsq7b7WK1ScWIg7kjulkuRc1LiLJT/93dAr67pOg9m5t7KRw++K1WzJFZHMRJANiBwBkhMCM6gjGjCAXhGDgIMwEB7CyhBYSREJgphljVNTPbQEoBACIzifBtsn0IYV+mDIkohGCmXddpyYAQY6WldClpUg6xbsZQj27eLv/zf/27X32xvu6gBdDvD/V/xBHfDwxq5X3MeWCT3a3v+81mIxJFBIEH2+fBmdnMeCdw1lJ2r4LEjIi+ey0cahYiAOjgxsM8rGp4J2ThkgshxhiK2uDdYWamCkPhQ9WHJUp2SXo7ETSAIxELx8gRLIBJABESITAkQhEerJjcrYqxripmBjdXlcAxSlUFc1MtOfewo8It59T3bd+auRsFi1siyeYhfHdv8kccccQR/8JwJKCPOOKII75xOHFSz8nNcpfRcglMo1HkUNXTaRyfjet6VNepT6UUcx9PJ7GuHEDMHJxYhCgihllxN2LiWDmAt63EKtQVorNqnBSIsxVsZqfLuqpo4JpvPReGym/gjCQcgkSRgIAIjMA5qzk4sDmhozs5gPmQjc5IDEQ+ZGKbw65UurAM2hcioqJqbkAMSIA0DHocMRdTK4AF3AE8pb6Ukksppu+WoNlv6QO8y0o8tuDXH0G8Z8mv0+BXUUnfzvPAjgMOLDseEtA76nk/jLzzfj4QMx/YfNytDu8o4gfU9P3tPNRS4t1W3TFwB1UM9xasPoxn3+nHe/JtfEiNDaeigYMI102jukYkBAe3bdsiIjMPNHiIQU3VTCgQkysOUiozSymFEFjEzAeDWiIa1sPMqmZuzFLXDSK+ff02q0XBqqrGs1nOue1avbqYzu382VP1UvI2t+vFYjE2CaGKk1lLctNdaco596IZQx1j9CI5tSlRVVWxDm232rbrkfr0SV2NRmUyUy2mlrqeQURiFm23W83lyeRsOp/Zaj3Kmz/6YPrpj5+l8ub1TfttpQB8VRBiXYWf/fSjv/yTjz98ftKur+sYppNpjJK6dr1eAkLVNCFwt15dX72GUFVN42CrxbWWFIQlVFrK4vVn7fIaShpPp/PzZxLo7duL9fKaCSYn89FssllcL5c3CjCZz5umfvP28urqMjI/ffacmbp266aj0Wg8nqxX2z4VDCHUFSGU1BWFyoFFzIwkuEcicfebxU0xbcaTZjxF8BgkxqilMzfV7E6q2cyIZKemB0AAZqIoq2WXC8M7OeH3P3x3gfc/E8BIZB5jQxwc2KwKXDMFxIAoiHUQJHBXIggsgaUKIQYiHMoDQBSKkWPgwCTCEiRIIGZ3BgBEDBJZBu2kDSrpWEURySkxcwhBVd2xqiI3FQG4FwQWrrghoFAwfHa5+vtPr//+s831NishoIC7u8Hvcmf6/nl0H3HEPxeG+9zuHuaqqlpCaKqqappmb341+GPQjp4G4UExQB4CAdyJoAfPDURyt8GXo6gaOO7lyHt6GiiEYTFmYqZhETdzMC2luJujvycE6+DZoctp23cjCA6qaBHQjdyISQgZfbc8moKCJwchIRQGIYiE1S6tIzgwDlkhiMQTJjQr4AAU6tOn0Mz+9ouLXksLAPDm2+mTI4444ojfZxwJ6COOOOKIbx4SQKiKUkUWKtpnJm7G4xCjBBGRpoqRue+6omoI9agJQWxfJdxhJ1sjdwczUxBR84IEhAjoaq7uQ60YAAkBaWCQ3Qbxy+BaAIPMhJhFJDBxTrnk4o4lD6a0CKiKNtRysT0dg4Bk7u6lqKqBOzMT0zBKMQd2KKqqpuZY1AGIyBzMQHVPDrq5GyFqKX1OavpuEiYAvIfr+Woc9HcCv5OucnhIOv8j4ff+u13r7c/3tuCAN/7ah2zPMe8l04/Iw79aO/sN8Z0jJYAjAqKZWzH1vm0BgVmIWc1KUVV1cCIOIWgpQ+atueWcJ5NJDBHBCIeTkQkHt0p2ADdDxKoZcdMsV5uu3VrqAtPp2ZPlYrFer1LqkWB+dsISYj1OfVquN9kWT58+r+sRoGzbrF2bcs/9NhBVdQg0Wa+0z71tlrPZPKtu2q7Lri5VM2pGEzBP221qt912O52esAgL99u15r6qYuw4eH4x5r/66Qdvb7qbTd/m7xAFjQAh8MvnZ3/1F3/48Q+f1ayd5cl8PhqPvOTNdrtt2/nZ89jU5tp3q+3m5ukPfhQit4vF9eXbEON0PBWWzWLxxW8/Lf12NJmcTOfVbNZvFml9k1M3bpr5bKpps1pepVKq8Xx+egau7XqZuq6ZzZvxuFsuuu06xtiMm34wKdp2zWQyns0ATFXdaeBKcp9KVi8GgBJCm9ZEHGMlITiYuYUYS44OkHNmxpx3HkeIxMKI7l4QTKKAOxGxyDuH5LvLQR8EnO6+DpcmA9REY5EKOSJGhshcCQeEyByYhJnI3YEJg3AUCcLCROhEIIIhcAxcRQnMIiwiLExI5oOfEsYoA/ssxENESoSJgAiIkAhUHdGZSZgQvCQnQuEYgyiEPsGnr68++e3FFzdp5VYQDcDhK5YG+M71xRFHfIdxF5JW1ZxLXcOeUN5Hu3d2Obvn0aB6BoChCOE+Wge3ltBDLtxg60z7lCz0XUDa3IdKpvuyf3uSm3h4HTVSN3TEg2jSPrsL3AEUvM9523ctmKEWMDVUJikkoiYCLi7E6Ag2UNCCTEiCzGiMJuRBQISJeQjqs0iMoaqilewAQFLPxjCevlouS6sA/xfA02++L4444ogjft9xJKCPOOKII75Z/PVf/3Xit+OYPnj5wcnJGPtnng2BMNbghuAw2D2XxDE6E1QVgqMZqYIquAOh5VRyDwBmmnOy1nLJbZeoFWLWXErJWnLxeLEsXddm1eKuuRgiEoLBPr0RkYhZBqpltVptt1szVYViZmolFxyKiftu0KKqqhpCAERVNVNwEBFiQkTVnU80ESGguae+R8JRMwIEVU0pIYKImKm7EVHOues7fcQE8NvH/+AWfO3F37fguzzXO3M+YJ8PtND359+TxOhwUGnQD9TVjzpB76e6O+635nAbdgLp/Xof2ZEvVacfmEE7mHkphQHAiiVHHMxnh/CGpNK1XTefjgEJmAjJCIWZCcHN3UejkTCRe11VJWcEYGaWUIqKiKuZmnOg0aiZXr+5vmpzmk2n0+lJKdq2675vu83i+uJtVY9CNeYq67pdrVYnp09q4tCMpqe2vNRcEnZbEg6xqscTNesX191qOY4xSuwo9dv1wr54cv68rseCsjFfXq83m02I9WQ6G1OT+0Xu1iwzRgoILPBHPzj/5PPF55frVzcb++e/CnYgptlk9Od//NN//Wd/8GRea9pOp+PxZIzEfWm7VAD57NlzkbDZ3Gw2yyri6enUrCxvrjar5Ycf/vD05MSJLxeL64sLszQ+PedmktXWF68wbRihqpsY4/LN59v1KkxPp6fPqtFoffEKUjuOcdyMStGL169ySqOTuVJ8/erVONRmjkhVrNQKEAmFwQui77rUJit9KRpDiDEqS0op51LMdjkWiA6oqimVnSLffTiFwAsYmGVhFxamOgTFh1cFHnz4znTVHrjTN/ohB00ADCCIASkQ1cI1QcUYiCrmKBJY0B0diAaiWUIQRhrMNwh3FtIEiHtuiogICRG1aM7Z3YYEeFWNdR0kMDoMdZsAACAASURBVJOZ5jxk7Jt5GQyB3D2X7GpWSpQwXKEKoe/1Hz5788mrN2v31qHfGcQeLTiOOOKfFA4Atrf2glJKSmn4sN1uEXngkFMpgLgry4FASEREhMNj2vbSZmF2dwDLpeyi0gNBPdwdABHBzIo+1DYPMyMiERjAQE/fAzrsahXSkDXVl7TtfQOuoAWtFEiMgYmJYwglxurONcgVzZ2HAhIwmH7gcDsDQAIw+P/Ze7MnSa4rze8s915fYsvKrAWFheCQINFNNocacUwzJulBJtPfLZPpQRqb6baZbjbZ3ewmtsJSVbnF6stdztHDdY+MKhRAAERhWmb+mSFREenh4e6x5L2/+53vIIxGbNScHJKi9x44gCoqAsBys329r8WkSZMmTZoA9KRJkya9bl0U68/7Bz8zz0pLFHw87FgIBENzGOGB+vYQu7auCiD0kppmH4O3lC1pGCVJiirJGA4hHPYHJEQkZFYFRbTWhr477HdoF7EjCT1LcgCJIIDGwdRynAAQm1xqjXVdrQRsrQkwiUoSkQSQebFqDgAhZubsiE4izEyIuffg0VeTjdmZAI79ZvLkpMQRVxpDRAgAXdft9/u+7VIIP/zL8aL+JFT6mg2+5oHfjVXl0vm3ABTgc4BXeWP1Jb58Cp1fAXnv7v0KKox32ZCnux8mlkdSfXqILz3X1xKj0Tf18kGNQdUIrnClmUm7lxiIcTavWu8JMfa+3e3LolBVQUxEh6bB6BHQMItAgsGgRYQ5czyGCIymsCK+Kqu269qmqS8UyvrgY1CjklqfbJKHD99AlOvr5973t1fPHz5+x7pyuTwnoKtnn/d9O8dVPVuwtcH3h/1OIUnqfS/EtS2qugo7H5998cXFo4fLxdL7GKLEvjlb3ItIqa9kNk8xEYF1XJRV7GcpxRR84dz52b1mvyMyf/mjR5/fNje7po2vXHL470DiqsK98+Yb//v//O9//PiisuLQPLh/YZibw74P0VWze6ZYnt9vNrfPnz3tdtfv//ynbl4+/+Lp4bCbLRaPHj92Vdm1PaHU9SwmN5uvSLFZ3+7Wt9G3rpwXZRli/OKLz4PAj958d7m61+62zz9/ipIWs3ltXXNz8/HHn7z70/e6aJ58fnl5efObX75fIQFg33siRWBrrWEmpOVyuS3Kgz/4vu+6brPedJstSELjYvT3Ls5vnj7Zbbf1clVVZUpSFAVJVGWV2LX76NvCFojq256IkmpOzn89V/eVL+h3J9o4xLcPIUunmJwQHVHBpjDGETk2lWULagktEwFoSsoIA2LKrQdzMUJuIghMSJydjYqoiECMbIiIiAtiTDFlAE2MhokNWWtCUFFiAwiAhNYYIiZCEEEAQxhCTEmj4M2++fDp+oOn6y82XY8qepcl/6+O8U+a9P934fidphBiDDHaws2Xi9W9s74LucWoIqiCqAwDCyJQTaowtBCUoQYqd5MeO0rkDg0KmkIiJkIMYYhpO5Wq6tgVmw2piow7fPE479K+ZBhVQkoaQBUkKQRBk5RAjE/Oh7wajaCWyBoqrXHWWEPMyExmvXfOWGesNUSABK4orTXGGsZM5bE0yXCISRT1F797sF32r+9FmDRp0qRJWROAnjRp0qTXqwL1/dXH4k3o+r7tutsrAyxR+74z1jJziqE57Hx7gNUSCbq+W29uQ+hLV1hrECGEICpIULoixtTs94Bora3n8+z1K5cLSn3qDo5LSOTbBlK0CESQJA//AQAQATFHNAMSMlNZlzNATihACqCq0QdVtdbl/uIiaq0tiiJ4n6GzKwoi6vs+xTgYnxEVIMaoqs5aJBKRtmkAgI3JcDCEUJbOGBaRpmlV1BD3/ypMhd+NQX/vh32sp5+/kJrxCn3lvO27POFL9yGofuXT4wv/PN3qy8z0Beyc56jHLTNoJ0TLxhhbcOF92zSHFHpnWEQkiaTETKBqrWUmUnDW9r7zXQtQMHPbtmTsUsUQxxhvb2/u3XsUQwwhCELXd6UtY4x92zkflIr/9s+fNYf23TcfvRP07ccXy9W5AKzXa0lhd3u5OLtvXVXP5svVot1vrlQWq/PZfLVY3YsCkAIhGEOq1HlRdrPlWby9bPa7+XJRF4U3gAi77aWzlg1GJSTXN81GUlm5qqovn191YV/P5rP5QlRTr2+dz9574+yjz6+e3Oy/cnXgB5RheuPh/f/4m1/96mfv2uQhJC7MYb8tnenaw6HpmN2bb//IaEzdHlJ0rnTljLzvt1sRPXv4hpmvMHTxsPFtA8a997OfL+7d732/2+5EkYw9W62I4Pr6uo/44NHjerVq/OHZ55/sdtsH5+fL+RIUb9a3i3vn20h/98eP/+4fP5zV5S/+gouyApS264LviNkY51xhmG82m5RSWdZVPSPDVV3ZtNjc3uz3+9lF2u93AMBsiJjZWEtX10/bzaaqZoygKTrnqmrmbAkobcOqhAAxhD/vs/2nPjov3PwevkbGN8pxTQcMYmFMaU1hjKUcmEoG1RBawwgCKrm2nnOWCYBIUgYYmDQwIQ9cWrMdmihnuTKRZaYYIxExE/FQyp/dj0SoQIjIRMYYY5iIQYQQnDXadCH6PsLzm+0/ffjkk6vtdRs8ouTeqSPY+oreAJMmTfr2OjYVVgVEEVHQsirni/lisQTYp5SMMUNzhfGjh3nLGBWRhsitY3CWAkDu0yCiSKg5O19BcczueHFh+m6dfFjxzkPRV46rMC+8MwAiMRtig4qgIAgJAQBIEUQhSIiKoCrJGnaGOx+tYWs5D5slReuMczaHBSGBcb0xhpmcNUSUEGfQsLeHPkbNPGSK4Jg0adKk164JQE+aNGnS69UcOgyz6NfNBtt+fbh5ToChD7vdfrlaVlXlfR/7TqPfoVhnkLEsXGFN6VxMIYQAkkBFBdBhXVWzetYcDoqwmM0ObQt9XzpnmRHAzc/3qb2+uW26Tsa8heN0XgdniQAoE7ExipAkhZBCUkR21hhDIhpCz5yNzyHGoKqZPiOA9x4RM30eKioBVISZQTXG6IrCWZucA4Bjpqq1FgDz5EQkJUnITETypVLNr9Br5XF/kgd9eYOXDuaVUPjr9/nSxnmzBPAhAIz25++AlU+skF8VknEaF30X5fFC9sAxMxwwZ0qfmJn15b28mFpw6sUckh8BxmL+7JrHYd8qkrzvUycpEWIaoicBEYiImV3hyrI0RKTiytK3B+ecdQ4AnCucc8RGcYyTPh4GESgaY401CCC9bwN8dNV88NGnT66b/+N/+qV8fnlxb1HNVj6k66dfpBBsURZFVdeVxLP1zdV+u0bAspwhW7alj6Hr+pqMYGJjrbOaiqbZ931Th9KUM2Q6tG172Czny7KczRdnIWgIh8N+k2J57/yiKKpd0zL78qyu6qrr9/cK/PH9+Xtvnl/tmy680g/2wzFoBFgtZj/78du/+av3H67m8XCNKaGSxBA0dG2jYKr5spotKLbr68v9fru6d4/q2eHmMvWtMZZsqUjr68vDZi0xLO5drB69lYL3XSsxsS0LWxtj2649tO387MG9t99lQ7urZ9vNtSvLxeocgPa7Xdv183uPfv/Z7f/9Xz/8hz9++oufvb3t4nkFICn4BCmp5HcQZPQpIgSa6zqcdUEVEdna3A0vhkBE1loAJULf+77vi6IMvk/RG1cwGx/i5uq57z0ZBgDzcgz0S9cpS7/i/lfe/JP3fzcdP953lSgIwACWqCpd6axjMowqqe8DW4NsrbUACUkMk+FcYQOgIlGAFdUQEBMxI97VKYwRHETGGDaGmWMMKUUiKgrXdp3vYkoJ8qGoWGuNsargfVINKgkkqYoIRWUv+unl+m//8OHzfdcDRkJIqpApFuJQDT9p0qTvQ0M5Wv7SJLbGOVdVtbM7GD7abK2VHGs1epdzlLO1VocFYxxL2TSnrjEzAKSUs6ChKDAXvpFzCq9YQxojOIAYVSSZ1ErK9XYnQsipPaAIkI9zUVdOE0tEEiJgBEtsiA0hgIKKSiqsddYqCBM6a6q6RNC+bYiJGUU1pZRCivu9qBCgcxYJo1J5SHYeekZT8u9/+eu3nzx5rS/FpEmTJk2CCUBPmjRp0mtXhBijMBACMVnLiAxILgk5B8ZYRldYlMQIgKiErrZMZK2lECgGGHvC2KKw1jEzupkiuLqKyGhsUdVI7GYLXtx/1t00UbxoAkj6Qo5DbnAOAEw4cIQkvQ9dFxQJUUUEAFJKXdc7Z51zKSURBfAiObhvcK7IWFCZHdD5USICCkmEmPq+R0TO3CFJEhncdoghBBiKOl8JWL+K7b5sq3mRBuMLeEhPth/8OKftbr5KXwJMLwRUfPnYvnwoX7FL1Rdvv3QLT7CuHy3C427xhUed2pB1OGuFk2twR4m/PiPkS3fheCC5ChaPnmw9OYIT29JXREWMBf0DfMYXX5nxNFWYDSL63kPsHIIrHIJIDPmtntc8iAhwbKapgMRFaVzhUkqL+Xw2X1hrUCIzW2usNcZaYiNJnCsBgNlYa31Im0N4vo+//3T9yXX7xuPHPzl3aOzF2WwxX97y8+D7ZrctXFnXs2q2aNq23W+79tA2W7KLsqok9L7ZEfeYsKhmrigkxqKcxb6NPkpKbA2ChK7pAQzZqp4nweagzf627zpJslrd63wM3nvvrXPO8szGt1bVX7zz8JPr3WfX286/nMQxXuMfgsY5yz96641f/+V7P3/3sYHEzATKAkbBN42E6Oq6ni+IOLTNYXMbYiwWC3But9n4rjNc2KICoK7dt4ctkD178IZZnB2ePukOO02xKOr5vPK+bZqGyDx48516ea/dPttePe0O28eP3qlmi83VzWa3I1d24P7rHz77m3988vz28PjttOt8TWJZ2FrDtu1EkogKgLrCphQVUi7WSJJU1RhDxgQf2LCOijGlmADAMCOAhL5vD2QsIPkY9/uDxEjWhBByl8t//dKXeo2OkRyWqbZm5jKAZiJEFQAFAmQCRlAAVAUhImtyBgcggLO2KKyzzIxMAHDsJYZEBAAxRhHhGEXGDySkru373iOiMxYQVSVFUQkSZaDWTJIXDmIELrzS8237ydX+48vm0IsAyl3bQQWY6PNRkw38W+kbXq7v8e31w79Tv+E5vrgZAiJp/hJQiD70fZ9ClKQAYNgkTDnfmRGV8h//nM51N/whxDzMy01c8/YAAHiS7kGngw8Y/tiPgzzCcUiDKgpKMhRYvKjTroQpJYkRRQyCpRwzDUzoCK1BY/JolJlsVbjSOVUhBGu4LJ1hwrlDVEBFGtJ9cvi1ZWbDgChAbnVG1fKm8xHgF7/73Xa5/GZXeNKkSZMmfXdNAHrSpEmTXq8UhU0UMmVVGhc5LdgUolAtAzKzYWvYICJo7H1MMYo454yxhtikJCLELCIpydiCHOs5ISGhFmxM7G01s87VxsHswt5IQBsAI0BUSEP1JOA4hcg+GCJSoN6Hpu0OXXCuANQYEwDEGNu2dc45F7JtebS5IBHlaI5xBjKEURNR3/UpJWbmnojQ+8BMxlBKKaYYQ2SkXMQNGWBLGjrevKyvnde9Cg7hMVtkuOJHyw8BAKgA0tCmXV+YnB2nS/iyjVdHfo0voddvBqcUj2fxMnC+w7rjb0+3zA+86/435i2+AKBHRzHqybENP+kU9urd7+AIjBHv0PELF+N4BY5mpbtfnZ4bjFPLF7zQd2dxvInDm25k0DruGQBEiqK0xmUbvbWOgUFiH4NISiJJJOdpdH1fxmjYdF2fOyMhEBJUVWWtI0BCtM6xYWOtLUo2LnlflqXv+yiKZJPirg3bTq4a/Xx9+D//5p/m/+uvZ1tfFe5itTi/eLC5vWkPO0JgfFjOVvPlPVANfbNdX8/P7HxxRipr77s+Ymyss4wlO1eWVerrFFPbHMoFzWdV4w/9YZ8SLi7Kh48e7jYqsWvbtm3bi4sHy+Vyu9vvdtvFclHXVQrpfObef+vi+T4cun+5jIf46naEr51BI8BqMf/V+z/9d7/46fnM+WY3c8YgMggnWW927IqqLI2zIfr182ep72ez2fzsLKW03x/aQzNf1cvlSkAZAVG4sIvzB8q2a5p2vzGIs9V5WRab9Y3vutnqwcUbj/u23d1cb26vfXeo6xpEd/td5/2980d/+GT917//6KNnN+SKJkEXUtt0du5msxmpHta3MaUMQ51zSSR/sH3wbdsCIjPHmHb73cX5BRGJSIwxRun7no0p64oJQWLfNGW9RCIFKMu62e+C933fS0rf+HK/9An6oaXHH6MQoGCeOVNbV1lriUgFEQ0ZMgyMQPlzm5PV2TKxQUJk5LKwZeGsQSYE0CRR85uPKMOjEKIMCbCAiM65GJP3rag66ww7AI2SVGKMKWFiNs45Y40OTXBRyfUBnlxuP748PN+Jh8HvOH7l5VL7SVnTlfhW+oaVRt+X8HV/LX9J34k+D/yZYOjZoX3XH3b7ru2CD5qy8QBjjDTEKY+FSoNBII8EUE6GB8PTDGMAQEJVyGM/Ikox3o0lhj4higPOzn/5B33Zf4DjUEMVBMCH4PsuFQYImQBBmMAosoIBcATIxIaqwlaFq5xBACYgRGepcrau5qBJQZCQDefgIENclgUAAKIguuUjKM70+bNNn9OfL7/NKzJp0qRJk76LJgA9adKkSa9XQqC24NSbonQp0nxhqxqJJSRgRsNHz536oIhiLSEhAEpOLBBQGUwpkiCTXwIkABRbGZXAiKKavGcbQNS4kkyOJgCAoU3V3XBfARF777e73Xaz3Ww2+85bVyJSSpKNzNmnfDgcsllONRe5EzMd5w+5eNMYoyIhxJRyx0LIUyBmxmyjExEVFUWAbKZLKfV9H1P6ZgBnNNICAA1AcwgipLw/AhroM2anDiAiEkISAQBDrKA5ljQ3S8y7xRw3CiqihANJz4/NyJcQczLC8RlzE8UM3wc0PGQ/4Mn8TAf8PHiIR6SMYxbji2R3fOhxWxzXCwAwPxFlvn5KqhFVge4A9HAUgIh6rJwf+86Pt05uHgM3hqkhwHjiw6bDu2WwQp2cW6ZXY2+iAZuPr9PdCwYAQDTU7g8xlENYBgBoDGF176yez8uqrjSxBo0JkQDRGGOLopzPyZkvPgHDBgGSiHHWWm5329B1RNh2/vpm+4j53mpeVbO6mqUQY4ySJPqgSMbZFGPXtjCfkXFJyQusm+6v/+nT9378bm3xbGbuzcs33nzH2mK7vkkxhL4v5ljNlhLjpu83221RnyHIbFarnLfNoWsP+80aRGbz1Ww2c6y3N5e77TpJvH9+AUW5bUNzONhq9+Zbj9vGsS2w77e7jajMlmcCcH193ffd+dk9Z3hWmrdt9b/9+4svbtZNH7ZN/8Mzpzxp/+m7b/7bv/jJWw/Out26IDTsWEFi7EMKIdqiqquqsHz1/Oknf/yjI7h///58sVjfbvb7PSLUs8o699mnnzbXV6Wjs/Pzal7vrq6eff5ZOmwe3H+wOLu329y2TYuAZV2p4cury8N2l6KAUllVbdcogqnqQ6TffvD042frXefntkgCSQQRnDGlczFEEel7732oNQFIWTiNHgCY2Xvv97u+aar54sGDB33f931fFMXZagUAdVW16xS6jkvXt01VFmVVsLUx9E3XFWVZzM6X7U5/aJL150hf+NQpIIAhsmQsIuf7VK01s8oZVGYUFGPIkLUGmClJYDFkmJklJq89OFbDlqmwRW4VYNghGlDG/G2huX8AV9VcVJE6RDTWsimMMQWg6Xtj2FqbRBCQmYGjUSUyvdLV9e73f3zy0RfPPUAaD3zSpEmvSQoAObcIAEBjDN73IcS+7/e7Xdv3okpMiITDX/78RzpbpgHGEVj+kdOzTgaTQ53ZCU3WO+/0mBo9jBByvxBNKklSSt8gfk0JIQ/dCAyxYTKEhJIDgXI2fQ62DiEMrbUZEVBUg/fMgISAKhJFgABzlZWCqIIgsfdko0FmpN//8nK5Kb6/Cz9p0qRJk16tCUBPmjRp0uuVIoUgFkmUk3IUhZiIAESAEBMkERXRlECEjGFrYwiaBJKoiKrwkEEgKAlVMxMGzGnOkkfzIaSQwPbYHg7DBOLLRzICaWYWFR+8Dz6lBKopRQAS0TwrYGYRFUknPWkUQETuutDkuUW+nUQAFTVHhQiAMlOKElPA0WZMQ6/CFELw3sur7c/wqlAHGD01OBp6EBGBONd4IxFkRzgRYb4TCSlKQgDLJu+DjTkaj0fyq6CaJNFg4x4pNA0U+jitEhVVZRpK04+k+o6E31WoHj2riHd4dqDURww9ZoTo6BEmvDO7jjAax9CTo7n77gIN74Ph4uoR++IdljqZE+roPtbRo3znvX6hmDafxLDgcZobMhinNS9miIpKzhfXu23uXrx88GMNPiFlO/mxi1Hs+7KqjDH5+VKMXdMedhuVGJNoShJ87L2xJgcpSIyg6qNHRGYSFUkpw/C+6zebdQi+mq0IQFPUjCOjTzHG3ifdRZ/yWkIQWDfx//nbf34w+4s3Fram68dvvVXUiyrG0HdN2+FuN1ssXVWbsk5t32zXhbGurJE5ivi+k+RBIiNaZ4vFwoc+bW5T2/hDWVZ1FJJD2+03V08/r+r6waPHbMzt9fPdbk3WiiozRt9DjNYam7Tw+qPz2a9/+qPrTbNvn6cfnEAbpnur+je//oufvPNgZsFEXM7nEGNOd9k3bQRTLZbOGn/Y7m6e7w67d995++zBQyG7v10nSXVdsuVmvwshNH2aLRb1YqGh3Vx9gZou7j949MYbkOJ2s266fr6Yz+c19JvQrDsf5udv/OjsrCjcZ0+fACja8g+fXv6/v/3D0/U+CACAiDRNgzUzQwje975r+6JAds7N5+H2VkStsWVZOeeMMXFMBMpZHK4oxPsQ07Ksur4lZmMtEqUUUorErIC9D866eV2itYRIxH/eFf3vAVQRUIEACMAQOzZ2WPYZ2gwSgWEiAsEERGzIWWYSQGUma40zFlUJQZUQmNgyM3GmUlaEVCEJimQATap4OIQkqe+9gAJ4os4YA4jBeyJiw5KXJJF675Mos22FnlxvP/j08vl673PO/QlCnxy/kya9Bo2JZAAAEGPMbTyctWVZNm0bQjDWIinmqDc4LjLDMQ/nuAQ9tCk+jjxOB4gimiN7jgvqp0Q7L9sTqgqoSJJXRKJlq8T4YEVIIl3wRkgJLaEhMkxMaFUFFEgoQRIUq2LYMFgBBURSQFUVA8ZgJtKAoIQExEqUV9EsW8MMTIYhewsmTZo0adIPoAlAT5o0adLrlQA6IC/JJ/Bem21L2OTRLjEjoYrGvk++JyLrXFG4ru9TiKgQg5cUC2c1hRg7Q4igkOOdVRQyA1Qfok8SFMuzfn2TkveaBOBFDnmEr0MH82wZRucc2jKJ5ErovCmNpDV3icETvnpafJrjN1SVDSOgqMQYVQURrLXeew1g7HCOzlpC9D7kflY4BGV8edz/intGJ3d21hAbY61FYhwANCKRMYayl4+zqRwzKTYZQCPmJlqGDYweaco91EWyA5qGROs7y2++nYaKUTGG8wU9Jkscs7BPL5CeAOQhsCSDFsRjdarKcZngxOV86lWiU2N1ZtYnSdKqkqH4cQY4zhvHTUZ0nhs/Dtue9OobI2TvAPIdChp2Nvwbx+s/TipBEFCGV3Dc49E/PWJtwNxJkHJTMwLA7JoWFZVIzIqoqpIk+SApGcNt0w/z25RSDKqSYhQVAIrBS98VTM65ECOC3js/L8siRd/3XgGGXBhruCzIsN95qdVYm3JIMBEgCUAv+i+fXf3dB0/vz0xpVu5ma52p5ksR3W42PgkbY6ydzVcqEPu22W8UAIzLZbwgKCl43xg756KeLc9Sin637poD29K4oowSvb969vmDN9+pytl84ffbdQi+79qqXjx8cP+w3QTfuWpWVxxiG/rd+29dfPjFxbP1dr3vfkgMh4izWfWrv/z5L3/+7vmiZE2ls5AEFMiwckEuFM4V9RxV+u26265dUcwuHriy7ra7w82tiJZ1XVWFJm9QhZhmS67qbrfe315WhVte3HeLZb/ZbDdrY4v52T1Xlumwje2OyCxWF6t7Z/vNVdc1aOqbJvy3Pzz5/Yefb5tONH9zKRtWAB8jxwiItrCuKAwzpBRjDDGUdeVsgUDWOHUFxGCtQcS+7/uuB0mSBBSsdXU9j5A0+q5tJSVEstY6aw8pBR8Nyem7/Dtczq/+1UtfdH9+rIqOfTxP7gAgAMvs2Fg0jICohphQY/TOOGZUSAqqBCbTdhTrbFmUhXM4LiZZW1hr84eOyahiiGMlSwIRIAKF1LY33vuQYpsdlTEBgIrElGIIMaVxJZD2h6b3AZR6MDddevJ0s+tSOPordehJOqU/T5r0/euFUQGGEL2P1trV2dmjN95o2jbGSOOiPlHuAQgiL3wkX6yjOtZPnfJnFAAYqsTwdANVyMaF4/gnD6A0D5FOMPQwlLi7A0OSbXMIiA7BYDZBm8I6a9gYUUzE4GxcVOWsZCa1RpxCUA6KTtmScWwsMjPmDivIhIaR1BgqXMn1PFmXGwP84ncPPn17+9pehkmTJk2aNGgC0JMmTZr02hUNGTHOGQOGZhXjmE7AjIiSUrCcvHHOMTMggoowGTaaHEgiAlCryaYUVaIKqbJqUk3MjMSFahSIQG65svvd7rDrvVcFJMAv+YwRkZgQgAiXyyWw7aOKAiITcYwRADLGBYDctsUYw8wZ6cYYRZSQFVREYohI5KwVFZEUYzKGmDmHNIhIkggAROiMJUQRORwO2+22bduUvqoP4alGEJqpjaCixoiiCJjgmIVBRMbQ4ImmI7rN9JYGtzMYZmM4O3Mx25wRVAWPSRmjX3u4SkhjjWdSlXwDcOioIyonvue7MAvFkyjnPGFTABxDpV9EXAOFGQ3Jx3rVE5qLqEdzkAKMMR16unXe1+CrzrvN/m0d8fM4GRzP8u6RozUaRtSfkbUeX507zzQc7VHj3nzL/gAAIABJREFU0w9R26cndXxNafSVD67yIZpbVSX6/WHf9b0iiGqSxIYLt/Btm0AJRFKIfRv6Lg2ZvBJ8H9vW1SWhJQQErerKMCdBVzjcU4xRQMlag2qLYqD7zpKdgTXHFkmisG76v/3j5xfL6v7FGd5uH91fVWXt+9CHm7jbzOezxfJsNptb4pvLL9qmUeJyvpzVJcmibQBUYvRJoo/JlFW9WIn3Xd9D01pXlmUZEdab3W69nq/uVa48W93b7XfRR65htVwa0qvLK6uxdIV31NzePF6d/+LHbzxb7377x0/DKwoDTj8j34HS3VnKXtqDs+bRg4v/5T/8u3ce368Kw4aKskp9bwyDJURTEBVE1pWxP3TbW/Xd6uy8XJylIO3zy7A/GLbVbO6MaTbbeNjNF8tycdaHePn5k9jtzy7ul3Xdx7jZrLu+u//ojcXyPCU9XF/5tqmXF3U9i1HW17fE5pDwj1/c/vU/fPj0ZtuHBACKCETVbAbcZxoKhNYZYlCJyffBex1bVuZ3duEsJodMMfiubfreO8PMBkSZTVXXPvVt6IP3khIpGjSE3Oxbo1hyVJEXr/a3vc7f8Lff5ypD/ixn+zMBGACDQKqkSIDWGM4Nt5CAGIlc5crCoiEUUZUE3IbU9I0mQQBmE9eHGIJoiinGGEVVJOVoJhGVpElAEsQYBQRIFUVUQpKUQAWYNbcNQELDbJ3xIcWEgPZ6f3i66zc++vE7Su8WRidNmvSahcdCLMjr8UVRxBitMWiGAV7+268ng4LjwAaGUrDhN3kIMNSRiSDZ7EKAY3UY3Fmgj8VXIklSElD5kgf6pF5sEBOVzhYoVgVVEFRT7EViYGNYICFpsJx63xpiBCYwDMYaa6y1JpddESsRGsbKWsOZkAszFWVd3zvw/GLbdiHpFMExadKkST+MJgA9adKkSa9ZqhKDISEVRnGGEDRbToYwDU2oQgiOGQljjJoSqBAqMAIRgIAigkljcz0ABWXViNYYaxnJAAowV5XA9mZ92/cdZgMLAggAnThNMj9FQETrnAuiJEhEZJht33uRxMy5hVVOpDgF0N77lBKTUdUkSVWZuChctuTGlJw1zCallCFwiB5AjTE8hgzGGI0xQyzDnwbQACcEOl/PBCmNNuPxpAhjGm08eGJJHhIzEFFUmSi7vymTUXqBxQ4+3pG6EmHOj8iPBVDCgWYP3DpncQAMk65xpqangc2qOL4OJ5T6FOlmc9DduQ5eoSP9PaZajBR+OIqTGeLx8PMDFI7dhO4mgHcRHAM0H/Z6nCaOuxgnoZKOjvfTox0fcOKpf8HzBHeTV4QcjAJ3AdjjE6TYtF3Xd8ayeiBmZ0zJvGOjmkglha49bL1v2SATxBglheC7aFkYNXiQtN1sjDN1WSyXq6urq+OcGJnLqqxnMwXtU8T7SyqsAMj4ZksAHzy7vffR1TvvvD131arrZ1VVzZZ1vfDdbeob8VVRGS5K64pDs03Nzjh7fnHhShMuQ3fYc/QphWa/L6qZKefFIh3aZ3F/mM1gNps5u9g3/X6zBtXF6uzhwzeZr2+urpvdobCGrVUG33czomXtbq77GYe/eveN233/0adP191XNCO8+yx8Kwb9siP+uAdEWC3n77/34//wm18tXSycKcvSFgWTImJSTQCmmpWFswztpuk2t1alvnfhyHWb/e7qxoqYs1VRz4P3t188ubndvvc//sfFfHX19NOPP/iXxw/vzxczlLS5vHl6+dwVxer83Fm3vb559vlTH8JFVRaGd9ut7325uPfpZffbD5/+7T9/Ml4ABEQ2XNS1sehK68qyOxy872IIs74FFYnBGBO87/p+TsaH4FQZQWJoDztQMUyFLUpXGuY+eAYEgBAjjpkVmlJ3aNtDu6pnoJBizNz7m34zfTt8+roYdEbPDOAQCyJHyKAEYJCtsZYBISpSVBQBTgpROh9ABEUbLyrqe685fImM7/q+a0WSD8EHD5pjniIqqh7DonIykCKpMYiMChgTAIA1CAAiAAjG5EgmA2SEik3bPl0fDgARCZFyb4OXzgVf+v8rLuLEqydN+rOkMixGZwztCgdIwyK3qGpOxzn9FA5I+bToKi9/IyKA5iaEiDg2rD6J6YAXFr6TkBAKYkgpwYvLrePi+ZF2E2DlXIViJKGkPLxAACLlPIIkMAgECpKycTuJggpIAjFJokgUFEQwTL5wTJSNE0jkimahVaVlLwLEALBd9a/tkk+aNGnSpEETgJ40adKk1yuJYgAixdAfIOzFH0KIKopIIcUYY4pRUyIFrTwAdKH3IYiqHRoJqsI4Uc9JzIpMDKBJ0Ck7NIgIxMimV93sD0+fPuu6hhnCXcrFMRcYEIaOe6rQdb73XoB4iLMgAMitCAHAGKMqKekxr1kVQvDHyUa+TzR2nbAhQACQlKJISpJyBgOoZldyiinFGGPsuj6EkPf7Da7fEfEMdHT4qTKkOhy5aPZTD6gTCccE5xNklwRR0mBwJuIBUw9W3+GkVIkoNyc02aIugjlKFYceiyNjHUnxnVX4+L+ROef5Up6G3YHnE0D94tmOKRk4MOMjrT6pS832pWGXR+w97lORTu3TI30+PsHgDB+Ac664PXFDZ7QOY5b3cCYvAeicGgIIhCfT1JMlgdGyDYo6zF2Hc82AmhCYiYl831sJdVk4w75tDvt9Wc2MKwQw9H5eL8qiVJAQe0Yty6IoS2SMXRQRjV4AomjXe+dcWZSmcIoqXeu9zxHUIBHag6R46vMGAJ/gnz+9/L/+5h/eOvsfrG4Ncl3X9+8/aLfYHg5d2y+XZxcPHy3PVgmi77v2sG2rsp4vl8vz6OOh2Zf1DNiqCBhXzhazZdhtrvu+q4rCFmVZFX3Xdc2+qquL+/cPh8YY0xwOSeP5g/O6mnWHQwh+NpuXldtsr2bVxU8erf7N4we//ehZ0K9F0N8FwL38LgMAZ807bz36zb/9y/uLwiRBST70lmFRu+awP7R9AlosV8vVKu5vQ9dqDAR6cX6OqrHrDKLEtFreS1H3N2vfdqtZXVibYkoplWX5xsOHpXOHtllvNoeu+9l7P5vN5uvb288++RiiX52trOH2cNjt9sp2J/a3H33yn3//0bN1I3KHyImH7Pne97LRzc0VSHKVY0aVNF/Mn2qKCopIxhSu3Fx/4Q/rerm6v1p1fdi5m5Ti4bAXVzJTDGG72Vw+e1aVVT1bZT/crK7PVqsYI4Uw1Cfot7rGr6hn+PYv0LfSmL8xPtkQvoE4Y6otl4YZkiHjDFtmYwjRJIXex853612jGkPv8zooqsaQfN9DbhablCl/eaacs1oUBTODkjGGmQjUITEzGwOgIpEIjGHr7JhrNNR5gA6RJmQr4SKgw11orjYBAIiQLUb/UgUMDjUY+Cev4YShJ036lhqrl0QlpeBD13W54o2MySljOvy5z/lsAOMg6jjYI5DTkcjxX3noCADMnON6xtK0Mc5rbJVhgFSMmJRiSCmeHh2MXxx5vCMpkaSZMXNWB4wgoAIIhi0by4aJkRkNQ2ltaQ2DECoSWGY2NKQ0pZhQsi3BMOc20t77JArERMxIopK5ednOX+8rMGnSpEmTJgA9adKkSa9bJMkrqYTDfkfdOhyu27YTAeuKY+KdJWI2ffAqEiQZa3MVIRDeuXMR2VgkUlXKv5LIrMwAY5O6Hio2nFJUUELgwdJypLgIqDlKObubQwh910cF68QkjZS6rs0O5RijqoYQRSSboAcUi8AZROQJjYhqDk1QBY0himFCCiFzhsFmHEJQER1mOTJmR3xDO+cJrB0hZ54d5YaEOjhwc8++3JAQB85+RL06WL8zDc0TEmLCu7JP5NERba0BgBhTviemlB3TR1ePjusBcGLzOU3PGImwZqMljB7nl36M3u5hKqfjnhFp9BeNm97x0yGrMW+AI2pGHVvPD9Ejwy90PK5jV0HEvN/Rfw16goGyvT4veMiAkAemf1eVi6ep1zCGc+P4Xj1pTJiXAo726uOBGARrTT49a22Ire987HsBYUY0HET2250rHBWlcZZ8f/A9I4IzZA32XdO1jx4+KM4WKYTeeyKTk6vzKy9JYgiFdQwAvqcQDEF+tXW88JtD+4cnz//LP33ifnZRuq1BPV8tDwTXV8+7Zn/A2+VytlguBfD68ulhuy1d4VxtjJvNlqhw2DdFjcKohFyU1WKx396ARE0hRXaGsHB9CJv1TVHXzrmyrNqmaZpuEaSqZskH7z1Se35x3vorhfh4Vf+793/y8fPbddN/vQv6zxci3L9/8Yv3f/pX7//Yxka7AxW2tK4qCFPTbq9SwHp5fn+1ZIm3tzeH/d5YtzyblfP5brtv2z2yzhaz+cX9ZrfbbZtD27/11gVLuPzso8vLZ4vlGVuHIJJ8koi2rB88SjFsby6b/frRw0dVNQPVrmsO+wOx/ccPnv3nv//gnz95FuWuHIAQHXPsmmg7LKqiLF1ZBt8Vxjk2KqIKxMyEiBhTtNaWZRkbAoCirJO0ufSbCDVJURZJuCjK+WKZs2EQUVOK3gcfEgoXM8yt+143QP4elT/xCgxQGDOvKmYWESUUkd57771ISjEkVVGNmkSSSEohWiZnGccvLkOGDSIpEzFlfKwIUDibV+aKojCGRQQBiMC5QjSF4A2Tsbl7rmVmVWVma8yxwMRU8ybRZzf7LkkASABRVPOP8TROSzm+/o8CAk70edKkby8ERGIGxK7rvA8xhBRTiJH6PuW+wsN2+X94rKQ6ouZjrsZ4e/wKGpbM4diaelyoHjZT1RzGBdlInZLqn/AfDLVbIkjA47COEHMzBmJgg8xkGJxBy8CITGQMWZP/KAg5h1SAGWriQJQQiYecEDJudn7PLJbxcMA+Pv7854fZs+/zek+aNGnSpFdpAtCTJk2a9HqlqE59G6P3Hvqub9u27VRJyVhrjbHEVDhXsPF9L0mMMdV8VpaFMWYYwedRPKG1lohVFa0FJpAIGkAjEKmIBGEsy7JwzgwJDbkRHt7N1/HO0Aq501sIPiQVhRgTALVdJyIlAADElHzwkpKCllgxUUwp73Ag2jpMWnJzq5RSCIGFiSiGwdvChkEhxshEOY0hp7Z+dYn711LpwaKjiKCYOTIoEYxEGZHuJio8YCYYbcU0zEOGDEQkyIa9geoOqBWNs4iYUsqW59ylEBFEZUjBGB4xoNXcukdEXgDQeW9DVelLtqEBhOopqR3tx3AaoXic+MlgHx7Zb95AToItYGzSOJLoo1n8znt8hO14mvpxSqAB80aKx+koDl0Ij6mNODLn0c6cT/VFMIRjFgnmjkZH8AsKahCIGABiEiAVicG3oe+MYbaWVIP3wYeymiGwiqokVXHVXBRSEiRSgCQxH0BKKSXxPqQQARCLAon6vqvK0hLHEEpmS0Qvvq9ClMv1/j/9/Qc/ur+oLZUMy3nlinI2W4IE0Ng023k5Z1MUxUxCbJuGt9uyms1mCwC8vHwqGW46J2pdWdZ1TeJD6GNK1jkRVe/btrm9vl4sVkVRlPWs991+f1guF1U979qmD3Fx79583h7aWDG+99b9n7/75j98/Pnm0L1WBF1V5Xs/efdXv3jvrYdnsr+0EueurgsDqd9vriH2la0XpS0NhcNOg2dm5+ari/vGUPTdbreWrrl/ceHKst03iFzU89W989A3+9tLDe3Fg8eKGGIIobfGvPX2O4bN+vLZYbu2jIvFHNl437dt14W0b/E//e7Dv//g85tde3xbIqhI6tuub1suqHDWOuuKIhIigCTxve9DjCkZ45AwpQSobJjYqKIkCSGyYQYmJpEYQyBEYwyRVZUYY4xBRHJWfVFY6xxSGNeWvt+QjO9Xdwd3/IZhBGe4risA9SmxsqQIKXnfh0yaRACBLOdgflIsncnZ9ExkjS0L54xBAEKgYbcCqM4aw0RERVEYY1JKoEoIzjlVCYasI2OIiKyzzJxSctaWZWnY5DIUM1tKEzbt833wGUAnlZR06EM2LsKdnN2kSZO+b+WyLyJE7HsfQ9AkKpJi9B6TSBpHHF8JoE84NMCQ14F05w94qZzqVCcAWnKOj7x6BPjCnaKaRERRFYBG3wSMVSrH1s6Qy9og+wQMIxOAqrPGOmsKi5RTOtLggzbExlhXFsszni17lSY2ffEEDvf+zGs8adKkSZP+pCYAPWnSpEmvV0okhmzQarZ0FeG8UiC21pU1GYOcg+yAFDRGRQAmMkxEYym45sSJzCdBEkqAGCEqJA8ScvZETJoUzLxazKqL8/OPn/kQQwIQOInrVVUAURVR733XdQjAbBJIjClEAcDee1FBoigJAPrepxTzo4goxpR5qiTJRlzDDAAh+IxfEbHpWxWp6zoz3LZpVRURbVUbNiGEFCXGr2k/+KcK4BVAEVQGb40g5vJOIBzuVATKGRCo2YWsmVoDZcCiI2UFEMwR2QCoioCoSDEEHKE/EhomAABVQwwjJkYEIj5uNVzdoYg189jR/6MnluCT/44MOt8x4uOT6d/dKY/kG0avNwyuwfzmUNWjExqATnZ/ZNw4zNfuAqdxvHs8chy3OmHVCKOHPL9vdAhhhPxDVXPje8xJ2TB4qO+OHwGBSE66EKkCkKa8YhBDFCfEiAgxBgUkZkwJQyJEZoOiqQ+h94xQFiUoSEwgQABd29b7vSF21h0AJEWVBIhgLNCRwgsmKVxBSC+95RSg6cM/fvzsd09uF8X5wuHs9nY2X87mM4LQNOvNZuO1tGU9X55ZY3ab9eb2xjDXs6VUMyTTtq111oSCgAybxdmq32/brgHpl9YBMbGJPuzXa2dcUZUr5n2z2+/X1nJdz5Rof2hVYLlcJtmELjxaVr/5yx+v94fOh9anr/sU/BlioscP7//6lz/7+b9527F2fb+YV4u6ZNTdZtNst/P5rKzq0hkNfbtZoyRXlLZw5dl57LvUHvq2TTGW9Vz6DoIvi7Iui2q5ury+1NAvquLsbNm37aFtQpTl2dn9R2/tttub589j8Ger5awuD03btV3Xp32Av39y81/+4eMnz2/DGL6R37YppsOh8T4xO2Nsft8TUZQUUiCV4H2KkcqCEFP0KVNNY4mN7zvve+IhLF1BmuYwKw2xAUAfIggkyYFEYKwpq9I6i0TfyV37A+Hqu6dRGheKhvsNkmUm5hjSIcYueZAEKaoky1zU81ztTpZVEqqWxhSGLKNIQgTDWBoqHPHQaFXzVyKB1JWz1gzfZpiUtCxcWTgAICbDC2ZiJmMoxhhjTIJF4crCDT1oRYJv9k1zubnadW0EkKG2QofyjfGsUHH43p40adL3rLHgSRVUmQnU5Eo7jgwAQEg6DD/uPoGUu18A3XWiyH/8Bx+0jq19AYbyo6EB81gHNWwPqunlb0h86Xvz+Ki7eilUxEQYkSNCUiVRRjWoJGkYxiUFRMsk48AQhoFLTgNCBFBJqgkBLGUO7SEhMTgGJqARtN/sHtX1/vu74JMmTZo06dWaAPSkSZMmvWYZ45VKp/ViVSQGzwBIxtiiBCLI0/2UNCZigwRoOKbovU8xiCSVJCnmfyCIStQYyDABaPKoCUEAMApExUKq6L1zjolVQe6AxUvHpDHGEAISWWvJQEyaAADIgYoIZe8wgLGGmAAgF6cTD4biYYyfPTV47CalRMREMrptYGSUiEjZnkycczkA/wzWoKqSYAjEzsHYBJI5KCFippsJj+kRw0woz0qyAxqJiBAARIRGozQiIQ0BiKNhiI6O8dF8jDmYgojghDOftA3E0bk+PPA0f3iIgb7zKEM274yb4xBVcecsOt318fmGkI8MoGF0bSIgoOAIso+pHGNUBhz92MdwkvxKDggIVPGYG35EyAD/H3tv2iVJcl0Hvs3MPfbMWrqrFzQwQIMERELkzOgczR/R/MjRn5ijc/RFEjUiuIgg2AQa6KW6lsyMzRcze+/NB/eIjKyluxrsAjDDuOdUVqaHL+Ye4R5m1+671wEIHEZV9K37BqD7wSxytLo+bgPHi45IJ59AB0Qrhkgs7AgSAmtRJjPbNc1svnJTcGVCEUJwLUVTdi0l5el8Ie55u+v37eWD+9B2XFWr1aptGhaRGADA+74Uvby8DCxt14fpwlHU8GVNsTrsEvznn//Tw+WfvXc5jTfXxHyxXPpkst9tn19f0SZ//0c/vri831X1erPt95s0ndSxYpaLywdXz79o2oaY6okVktlymXJutjtyp307mS2qSkra9c1+d3Nz/4MPJ6sVbajrbq5vnnEMUk05+27XLJYLIqDtDtr0Fz9857Ovnqx3zZfPt29ikf5tQYR1FX72bz7+X//8x+9czpr1janOFosYqNtv9uurEONkvqjilMm1b7bXz7QoVZXUc5sud7/6p+bmupI4vfeQ6un+qy/b/Q7I43ShUvWpj4zz+TRE2V23T58+v3j47rsffE/Vnjz+crffzabTBw/eqWN89uRJ06W28JNt+b//n3/8x98+2zZp/HgcuRJAd0QOSS2lzBJMCzL1Jc8IZ8tFyirMgYnBSu7VTAG5noZJXTQLQ597cKhmizqG3XZbRQxVXU9n690+TkKYVBxYS66ryh20KLiONqFvit+fTPpk1misIxgcWhGAERkBzayoq0LRokbuBEjEyMxMwhEJiWmwZqoQA4EQEAVEIPQqUBSKQRCdEIIwEwhjHQMzA8AhIaBUVajrCABMFIKMLiiEJWNmKEWjYGToSzZVAEip3zbN1Wa3T6kAGJ6cEA4zcIc5uDPOOOMtwQHcTIuphhAIaYi48JOvawBAv/vn7a/DPgZbIz/+fmrHcSCd4eQZPq55OxkPd/d4p4F+7HUM02vFvOkTGxmREDICE5orDyko4I7miqJGaG6ubmquboFJCMy9qFJhYmRCRxImZhytQEb1d0o5G5Tl5T7lP96ylzPOOOOM/9/gTECfccYZZ7xdOGAUqrCazOcxe/FUipq6lWJjUJtrzp4P4UyEbdt0fZv7VErWknPuVbNpGXLIzXUwuXNTAmdEDqIO2ajSyX67H/S+AIB0mj53bBEiopmpKiCGIIGkmJujI4YYhsjBgTmUEIYN/OAlPMhdx8Qah0FnwgQHt2gkZnAfOAtmDiHAQPIiDktkMB5B/p2Vg+7mhjAYUCAeotTpYA6BxzYfz/h4RkjkNsq3B0plsAdBIjMjJCIyt6Nfx1HMPB4DR2vpE43z6IgBB5b3dvlhwDXGLR4GXbcio6M9Co5/jYohd0A6Etjjj5FBP7aKYHBUPLitHA9OCESHlh0F2YfthyYNGfJwEA3BYcjnQwihO4xNQzz4pbg52OjtCIPNto9n7m4Hhf3wBt1+1o58/ImFNIgwIrjZZDJB2jfb/Xa97VOJVT2ZzhAgd61pnk0nRBRitLp6/ny35U1YrZiImO/fu5dScgRi7rteVVkEkAAI1UMI2+2GInGorZ5tmy/6lOxVoZcG8Pmzzc//+fGj1WT5g1UupU99NZms7j3YdEndNfelZGSZTGeo/XZ305dcz1cP3nmw725y6lJOdT2ZzSbIEmfLWbG03/W5SCnCoa6r0ne73V7Wm/nl5aSezGZzs3XWRFBLkN1+FzthxknNuWRB/8uPP3x6vXu+3nXlux8P1zF89P47f/nTH/3g0eVcYGd5tZzHwKZFTSVUs/myFBAuBLbb71O3D7GaTidVrNqnz7/4zW+95MsH79x/7wNEvHnyxebqqpovpovZl4+/3Gw3NWPNVLbrbr9FhJLz7maN4JraGMJyvqrryc3V1XazzlQ92/lf/9MX/+1vP9ns+5P3ZizZQABkqqaVe7/erNuuDUREVNeTup4AYFXXVVWDA4rMLi92jx/3Jbs6F+vaVs3MXViQqJSyuriAkm422+v1WmIIElCNAaqq2u12q8XSAcyOd8MfFrf3z+lSvPPa8f4EHpTDZtonMEf3YbpPCAOBIAB4DDIQxTFKIIKcBDww1JOKCcCUCYJQHZkImLCuYhWlCsxEiGDuMQRE7PteAsfIYzE/DZOS6O7IxCgZPBAKWJOTmmGQLqdt093s+jZpGR84iC849pzZ5zPOeIsYv8HVfDDJUWJmHsudhmqEk/7J+P+x3zPMurvbMVPi8HV/8qU/2mIchNR3cGLdfpLa/CKOtDUAgAGkYpum9UCFqeIgRMKggQJ4ADJwBTdHRHNXBiMExixCQSgKD5UcHChEERFyiCFMJhU5mWLfZ5A+Wbdv2tyrzvaVTf/F1/mMM84444xvwJmAPuOMM854yzA3z1BHJMDBnw7Z1DynXFLKqet7TclyGYLl1LVt9qolhkiMAOZWokicTogZwM0LEw9Wx4ElCLsPVhMM9b3qibqxOugJD0jEPqT/wTCsIDcvpeS+b3MxJEdyx2FwMqRIDfEvAINSmIZMQkIamMSRoiWCAsQEwoOoWN2YBpkzupsNxhwHBnUYeqhqKcXd4NXs88sLX+ImjoJiR6Ajg3uwnLiV5+LpLsbRj+rQEDycIIz2zQ7uCm6mg65Q8TAow7sNwNHkYmR3DyMrPPBBJ3T3iT75zg5OREInGvVxw4OO+qhIgsOCw8YIAEAERCdML56Q5mMp+6GBeKsxPP5/SGocD+/jRfODC8e48iB38oNttzuejB39VIB9Z7Lj8KYMF4YOp3g4MoM376xUlZi0qBvGENHputkMPuMAnnPvYGYFoGgpfUrz+zXXtZYy0M3ZAZgNIeeeCIgJ3UGLmyNSSn1gAde837gWPBlNv4Au6y8+ffJwMXl0bzHBnqzAYlHN5u99+L1nTx9fXz9R19XFvYfvvnNFpdlvm3ZniMvL1b2H71xdPW+7lva72XyRNVOI84v7ZTLr9ru27+po0/lsPptfXa+7Zu9ok2l9/95DcC85J98yh+mkapo9B6wC37tY7Hv80QcPP7vaP77Zf/LZ0++WgWaiy9Xy3/3FT3/4wYMpQ0R/uJpXkEq37Uoh5Pv335UgqW28pFKsbzYcKNahqqOgrZ8/yzlNp7OPxIhJAAAgAElEQVTp/Qe4XF19+uuu66oqLi5W9epifXWVu366nDLzbrtFxHcfvefI6+srTV1qm9l0Np3NzWC7awqGbZFPvrz6b3//q6tdl19Sp+PIjJhrsdJTpCrWMUi3vSop5b5PfU+DfF7I3XLqRaSuJ85lMpnMFsvdbm/mXHFdBzONIsBY1XU1mfSpV1NXIwAhqmPFg42+2eFe+aPF7YcYwcf6E/c6xmmIEZF4oJ4J3Qg8MgoBAxIYOVRBxJVNGa0KNAkigoPmOzDGKJOqQjQErwIFBkGvggxKSWFGwkkQACem2XSqqk3TALE5lFLMFQlnVV3FKEym3jt4VbXPNjdN3mdINlpCnRSEDF8LCHCMJPvmj/w5hPCMl/AmN+0b3thvuNobfgj/SJ4mRyaZmFmCICnLENlHJHI0rTpRQNMQeQ0j/zwUnqmPzPS4xP2WmB7+sKFDBeN2JWdVJTzuxNzV1caUQoe7XaRx5n7o4gAycihampx6T8IUGUVYhJmZCYiRCaJQZCL0QSIdhIJwkKHYzYkQEYkpSkQkB3MtwjxdLGYPpFpJKclAp80qYfN7ez/OOOOMM/7V4kxAn3HGGWe8XWjO7pKw2d7chHRjzY2rurq7Z81Zs6p6UTCHITnFjdA48GQSWZgASoxBpKoiiuAgUD24KwQWZjE1c3CkwlEL7HddzicGsgc3iFsXBxqUsN6n1PW9IjqyO5rBQMUS8eDgCYDExMwDAY04UIng7geHPSAiVXF3Nzc3ZiayoZ2qOoqBHQho2LyUMtDcr7lgr1z+NaM4fO06p7YPo5PErUWEnwytThtzquT9mj3inddv1z94XuBx6fjzTkEr3rbpdOfHAtbjSgMN7MfC1NvsQEcCpANvPZLJLxDQBAcZ04my89ZJZOCgxxbibTsPzhm3NODgo+KH8xilT+DmdqzIfeli4UgtoZ+8RQcC2krKg4NI3/VuHiQyCFFDyGauWgDMwQwUzMwNCKSqSFhT6lLat029WpIEZCJCM9VSTNXNhhaXXKxScIXST+pYxcBMLzYRAADU4fHN7u8+ffrBw4uLH99jTwY4v4j3Hzzc7W42mzWsryWG1eqins3VLXWdlq7draeLVdunlFLbNtvN2rCWehrrSYhV23V92qDrbDJdXlxum3bbbLP2RMuLi4v5fLm+ue6bXYx1CHXT7M29queL+SI9265q/tEHDz97uvns8fO+fJdhhLPp5KP3H/3FTz++nAX2XEu1mM1192y326jzbHk5X6009RgEPZeczEo9m05n88CQm023uQ5VmK+W9XRSUv/Vl18I5MvVvI5hf3OlXRtE6nqiiNfrzXK1Wl2s2rbfXF03201gWSyXsYpt215vtxpmn191P//Vk198+lV+1cPAARCRmREcTEOI0/kM3U1di5acc0ruqGbFoKiBO4sgogSJVRwmmIjFzLu2MwUhnk4rCewAJRdmKZpLzmZKRA5OeGt1+seJwxNjLIzAQy0FAkSWSqQavI0QmZCACFzI5SCRFoLIyAAMFgQmQnVkkSEbjKJQFWVSh8GCo4pDEAFGJhFmYmIiJqa6aHG3SYyllEzELO7gRd0BzUENio5fB4DZ8HrfXW2brljxwVbl1Wd2nKY844xvj+/2zv3GvfmbfVb/2J4nR+LYiDCGcKhLo+P5DBZgx8n1wxPnoGqm4Tv01GAN3IGOBDSAqroDD95l7kYGDnwo6DIfHdvMDszzyYX04/Q8gAMCEouwIxsxuBAxETMTMZIgOeLgJE+ANPR4kJGYkYe0wsHGyR3AjbKhu+VcNCcizBC83pcQS8oO1msCDL+Xd+GMM8444181zgT0GWecccbbhWtx6zfX3edph83Tsn1eUkbAGCtkkCiL+UKiEFKMQQKTMCIyi8SIMCjDDGAQiyAgIaKZmmrJGZ1MURWKarGcud9u98+eXaWuZ0Q96FdgHPYjgiMCIYkIM6WU2q5TRHMYjRUcETBbUlUzG40qmNxs2MFQrcnMVm4p3KNHx1Fk6q7HVwlxIKAJCYlSSmp2mzTzxjhVsB5C9/AwIgIYdbZHvS8ca0VPNDYnjOuxHvTlt+xYVQrDMMjvDCRf3OSEXz1WrMIt2+0jV3T70lHZfLLXUSB+Kr88cfMY7Eb8IDJ2B3AkAwIAH202DmzUwfGCTwxDwA9q5UMrBgn9US1+tK8ePmJDdf3ttfMxu/Cgqh75ewM/xAsOp3YQhh/+ONpDw4kE63CmAIBFlUpBNVQAg7qqq6oGRHcLMVJgZEZ0FgoxGJibgls2Xe+203uXzDTYvJRS1LtSymg5DTAEGyKCVGEym8QoX0Mvdtk+fXLzX/7htz98dxkJ1Pccq3v3LuaLRZ+6XNJ2syaEUE/mxA1t+na3uXl+f7qYT+fad836an19LXE+QY6xZolq6IA557bb1/VkKDlIufR9yHkym073u22z35vaJEQJsWh288BCbpDbd5eTH3/4zt/8Yvb4evddUdDM9PD+5U9+/IMff/TeRLpIXldSid90u36/q+fLqhK1nPuGcXwYcKxmi1VV12W/b54/zd1+tljNLy8ZfP/ky/XzJw/fuT9dLL3kp5/+ysxWF6vJfNH33bZLDz9cmJbSd16yO967/3A2m7uVXbPb7hudzv/+N89//skXT9fd684PiUIQYQYklhCruqQeEIiIhJGwJM25EDASSYjYJVVDsJKTllJSChzcbL9r0AkdhC3nPvVtSX2YBdXSdk3ftuYObszEwu6/g/P2d06b4oHhOnniwfH5Pa4BAG5G4AExIAXiKIzuaO5amCkwoRc0B4QYJEaphAhcgCqGIYQwCAkTIdRRqkqqyCIchOsYiBAdVJXAWZAQhbmuJzmnnDM4ENKknsRYgYMQpZJSTvvdvkNg4n0uDdCe85fPrp7ebLKZncgrzzjjjD8I3L3vUxVjXdfmrqoBQFXVFMb+yfhV71hGMvouENHcYOxi3ZlSwkOvZUguVbUhauNIQA8KaS+lbZusLwTtOoA7jgnSQ39SRKahmgpVTIFIcJQ/ExGCETqRx8BRmBGEUQSjDNklONLTPB5ah/I2dc3J3ThSTo3vMBkoUoGKIb3VK3/GGWeccQacCegzzjjjjLcNAgeCqo4PL6Zc9RqLFkNH5lCsAOEkRoDBBaKYuauxiFrWroA7IYYYEEHVihogMg+PbiRiMHd3EUICVOQqTmeT2XwWpAHo4Sj1HVMCR9KXCOu6XiyWi8VCEZOqxAqRtFhJ2Q1iXQ8ZeDllB0ckGthpgMF9mVnMtKgOtZcAACfZXYfyScDBgMTdzRFgUOWNhCi+oYbom3BLnd4uGinPl5mtsa3fdNyTXJ1xd/6aFcbjvbj8hGc5WB8fJESnW7601xPKCccSVTguGnY+GGM4ONqBkD5KnPHYGBw1pEOWIR5EyAhjHCCa2jEO7LQlPrL6OHwAcGS7xzM48uEntioHWdW46m27/cChw0GwfxBVoSANBpSpLxf1RLXruyb12V058HQ2VbAm51jVsaohJ6YQWfq2m7ZtLTJfzfNvTQ9FvwaD8MrcHYmponoymS/mUQSYZDbr842+ygD69PTXTf+Pnz/7uy83tUx/wKxpt988ffDOw6S2325L3z/76ukHP/pY4iT1ab+5Kbn0u2ZxcREu7z9tm912Sx489jDJcTJdLFeeWyx92+5vrp6tLi4uL2ddzim3fd9crC7rutpuqUuldqwmU+/2+31bynNCIm3n6B9dzv784+/f/I9f7PvvJhppPql/+L33//KnP/7g4coSLuaTGHC/W3/1+ZezSTWrK/Zy9eSL0u5FJE4mEqtqMZ3ML3Kz21xdb66vAPHi3r3J5eX++urJbz4R69/98L3Fg/vXT77cbZ5OYn3vwY9c4rrtebGa3n9485tfb549A5CHj95/+OFHzfb5+uZ6v9+ixF8/2fz3//npL3/zlb66EmKwbgEEIoxENUBwQ0cGwlDH2WIxXS1324aJp5PZtJqBghWfz6bb6+ftbrtcLl0NHOp6Mp/NtS+Bud3t2nbNpFWQSVUzctd12926rqtJXaGEoUzkd6JIT+6Kt4jjs+T28UKIkWjIIeSxwgDcBr0yoRGhC4IIBSYmCoyBIJAHoSpwjDJInUcmmnwgcRyUMAwO/giAhH2fcs7DXKOqrtdrGJIJHdS0aVs1NTckNDMtxZHUsO3Lettv9r3aK6/OKZ1+xhlnvG0gAJhpzrnv+5KzFjU1NRu+InGcaUYHNLw1mgcYZMs2TB4PXUI4FDkdd42IZjak/yGgjmEhXsAOempzVVN9ZSTDoYt07DC5EEbmiikSMgC7sqEQykA3MwWhwDRYCQXBKFyFMWOCGTmgRGEmYhr0E2AAru4GYFJFqiaN+tNt15Ycjf+v//Af/s//+B/f/rtwxhlnnPGvF2cC+owzzjjj7YIIEapZpavFMsTOQgEFcCLipEXBQwhqWrQwExKN+XHgJScAZCYBAQdXVVWHQYM8iFdRTU2VmdzN3BBBmKoYhwzAo8+m+8noH3GobY8xTiaTXpVVY1UjshfrqHPzuq5DCIjYNM0wThARJHIA1WJmIuLuRVVLGUjd4Yh2m7bnhESEpRQ1NXMeVIsIOWd8tRfCN+CosD7xy3iBOD38+uKrt3t4ea+vPNJrWgAAR6b1FHjkhk7bc7LNacD7a4rN/bjecQd4VLDDyfJbCfKt3hzw4HThcNT7OCCgDYz1QAUPYnQAsIPI6HbwOIQIDXsdiObjsPMwCsWDqzScjDlHM4+DkcdANB9F2YRgeDSydoCD0QERhRCm09raXcnFTYMgUpVTKlXUom3bgTOypLbZ7Xb7/e5itsRYOSET3btc9alLhHWsiKWqKpaKETX1wIJmuUvOmgHCcrHrupTy611fAADU/HrX/ee//uW7qz+7vwhhu22azaPv/2i1WjHQ5vpGc7l+9ny5Wk1nUyur/WazWV+beQwyW65yUS1le3OjjmEyn81nXi5K33S79X6/ni8m89kFEu/2zX7XCAmRTOdL6nMptlwuAlOz2/RtJ9V0NonW5AdT+vd/9vEvf/P4s2c3fS5f0/I3gRB+/P0P//InP/zhexcRy8WDe5NJlft+t92hyOX9h8yU2j2Dch0JsU8pO60uFiXn9Xq7bzuUWE1rDqHb3OyvnmrpZ7NaRDRnMJvN5zFEruo25bqu33nv3bzdra+ep7adzS6ncUJFc9vs99t9n3K8/C9/9ze//OzZvv+6mMXhpVhV0wrM7OZmDa5d34tI1/UyLdlKn1Pbcdt1Vk2bpkm7DYFPpzUzM8liRlVdV7FqkolwnMyASrPfZSvoQIQsDIjrzeb+/e8rh1LKtyvKGPH7409fdEsFEMTIxAQIju40ctDEiISOSEIQGAKLEDNiYI6CgSwGjlFikCBERGFgcwLFQCJUSjEihDBMFA2MVSkFDhxT27ZEVFWVqZZSuq4FBCRiIS1eskIIBtgn3Xdl3xV1eEn+fOadzzjj9w83MwUtWuwYHQgwVA7hyW15+jAcVhss2hyRboME7zwyj4VmboMN0sHCy2yYqHZXNzO1134d35nvH+htJwd0G/OQ3QAYkIlIgAOSoAu4AEXEyBgZhRDAhEGYgqAEEiYURkBwY4qEblY4MApyoZut7ry817//NOy/wwt9xhlnnHHGyzgT0GecccYZbxmIyEWd/eCAgEhEIhJlOnUmPMQyAREQAg+Z3iosRETMyAxm5IBMZq46SF+RiXJOqW+JKJfc9YV63m03fdeZKjqOStyj/fOoSAUk6FO/bxpzDyFwjObISGFSxxDcnVlEZOAxSymIGGMgYnPvuq5oERFmBsScM7gTUV3XiNh13WAOmHJPREEklzLE+kWJhKyqpWjbNIgv1pi/CW4HLS9yweigL/HNr97HtzriyRZ3D323WS/tfLj4/qrVDnLiV+4QjywyHD8Xd9bDw3gPCe/E9/iB5cbjZRqdLsZ/iGDodOCMYVx3pM4Hcv9weDPHF+Xi4yndGmwcWnzY27D2Me0Pb8np20YPkx8GXkoBNwmBExmTEWkpJechUC71PSIO4UYiEmNwh6qKDK455ZyIiYVJBo8ONDNGIKJhmsTdiZCIQBV2+0ldj1Myr4cDdFk/+fzq7z69enf53uJ+Zf3m5vr5w3ceLRbz0pftZpuaJsVQ13EyW+yatutaQqblcr64rKrZ8ydP97vWd7vJbhfqannvgeaOCPab667tYpVjNVnMY9+1u10bqnq+uJCY1pttyQnBmKkUG1LhVLNa+YDiv/2T73U5P77a6L/AiIMJH9y7+Nmf/uCnP3y0mkDfrMNFTWZ926dcVg/frRbzknrTUsXKTNUdhpRRxOsnT/quRYmT2ezi4QNhvH7+ZL2+AuF79y6rIFdPnlw9eYJcPXj0geXkfV+Bx5K//OLzZr+vpJotV5Plcv382dPHn7clJZz+/NfP/+oXnz9+vv0mdxF3d0ISDmi95RwCV6EGx67vqeuL2vDMHDztmajk7DkJT+NkVrK2262DTetqNpuYqqlrVu2L9rn0PbNU02nYb9u27bquYOm67utnKf5QGGeCxvki9IMBNAMIUwhCAGCm7kjExCKMrq7KRFGkjhKG2T83QhJiYYxBqhhCGMvVA3MMHCPHwACQUt/3aqpBojuklFJKqpr6Hg9OrCEEEe7aLqU0eD4zQpAIDikbSUCiknLn1Bn8Ds4mZ5xxxneNkRMmpqqqqqrqcyKiKCMhcOyY+Evz7O4O8VgLRXg7oY6Ds8YYW43jHJU7iNBoGHaYLndXM3PRvjV70YLjFW0tRRNAx8UIAqIAmGZVtCKWUYWycBAKQpHJlUELWTBCAC0ZOGHf42CNz0EAwEzrSkIY+qloxI1yLhkL/P3s6bL5ncQRZ5xxxhlnvDHOBPQZZ5xxxtuFAXgBqxFjzTwnNKSASAiEUYAISgKzkQYkApaUGu2TaRqsm1VNS9GSEUeD3tHS18w0mxUicIAgVLyUnFLfWSl4tI5wOGUpEYCQwMHMVBUAmFlTMQBgP1RojvmBQ8XlUHPtRxyI4DGGcMgKO5COA+UYMQIAIIiwOwM4ASFgCCGEwCII30VH/1Zn/DJt9Gpq+xsJ768VP7/5pocx3OuOd4wTfAVrji8tP5VWjyM5vA0kdDi9EncuydETxAd1MqoDIRKijyrnU178aJ490tkvOI0MFPQpK+3gt+Yfx5VGDTQc9dGnmipEI3WCkksp6gDELCFACQiwa1omBnMtB8EyEYvEEGOMROSps5xUCyLGELBo6fqScykFOTshMpVc+pSIWUTIHVKqwmsTCE+h5psm/c0nX3z0cP7o4p2LOE1937dNXS3m81Xb9Jpyt98hTCmExcX9m+fPU9/lVE9m89XF5Xa93e3b1Pe77Wbii+VqJURltlxe3N9vtttdcxFmi/mSUdbbrVOoJlWIKNLsthsmIMC6rkMMuZTAHqmfYfnffvzhs+vNvu3X++53Y0YJsarixz/44Cc//OB77yzmlZOba0655JQlVMvLeSp93ycy4wlziFqKMAhxu9v2XePuoZ7U82U1Xe6vH+83Nyl1VVVfvvuICXc3N7vt/t69e9PFxfNnT8F0EmN/c91cXzPybHUxXS6sdE8f//bm+krj9Elv/+mv/+mfH1/t+/w1zR7KwJGQmXNuBbSOkQlFBJHMwRyIRSSICAsH4UAI7qUUc6jqWS67tm3Riy3nxBGQCJ1BhIJrNzymSIhF1Gy33UE1cXe1V1tFvL6ZbwXD3fNynQXcnRASxIp5EmNAIgByh4EDIiAAQhz8ncGUmANT4BCFg/Ck4iqwMA2iQkJyt1IMQcEIAEpOCERIWjo3NzNEJCI7lM8TkZp67+aGRAxehRirEGLl0FE2qWvovUldq55eMjE644wzfv9wB3ezohhh6IxJEBY5Lb26NdwYFxyMck58zg6uW3Asd8JDz8TMiiqO+SFDCKDdPrcQCcnpVc/OQ4HboJtQ92yeiyUEBlB1JQpEDDiafBmCDh7Uh1xuckJHNBES5uE1NrRht0TEQ9CJOLDTMC3OZmgZUiHYbTfxTIycccYZZ7xdnJ+zZ5xxxhlvF2oIyFldkU2mUKmJuIGnjE4AiOqgBuagBkwQcb9rc7sD7d1NTXPOKaWcMzNLCCFGADTVnHIQDEIGzkFiqA3ctWhObjoEiaENlCGdeEQgIxKhIxQtRY2ISi4Dt62H0kgiQsRSypBGqKpE6O5lULa4uzsRlayISGiDCK7krERMJEKqmrUMTqSIWHIBhxAi3vo7fBf0zW0d6DfvDe9Id1/cxb+wHa+kwP3ovHFwcL494msP+03tcR+S/fDu9MLg1nEsiL0dUB4v0ZgZhG7DJMQQa3lCNONBAe1wa+pxaPbxA3T8bfRghoNu6va9OL4feGfHAACoiM5YStFS7FDUf1AotyzCwgiopTALimju1DSI9KmXPpI7EQkLI3mfcrHBXsPNHNwRVS2lNBQVAxFWVS7FXxWm9DIM4JPPvvqbX60+eufi4sMLkrRdb3Ae6sl8Nl9sd1dtsytWpovVg4fvdPumpNy1LdFGSDhEqeqctWtaQBIiYRau7j94b7/vm6afzNLFvaqazNb7tuuzeUvMl6uLJ0++ArfpZFrXE0BC8KEWInr+k/cuv/jBo+fr3a7tf7c0whDkweXyZz/5+PuPLu/NwuUsxBg096lXRJrP5yHE5zdXpW0nITpKNV+Uric3S+nm+fO6rgAwxGmQsLu6efrV49x3MVbT+WIym+f91rVMJtV8sWy6/vrmZhIkIvRdQ+rz2WKxWrHg9ee/unn2hXK4bv2vf/3Vf/m7X2279I2SWCKMIbBQu28nAWNVaUmllJHmrGpTFWIEQHQmQnAJwTWyhBBYtYCbuXapU+1Xi2UQdp3NZ4vdzT7GiOiqxcBDCH1KdTUJIZi+VEjxh8GxaODw97DkIFBEBwIISBWHKsRgNhShgxmaoiMzBuLALAQITgCRaVJXTBCYqhCDIKGbqoILU9GibpqxMCJCSYVFzDyn5ObMzCJMVACOk5GlqFtmERF2x+m0ruoKkFIuKBrqqZW03ndN0TxMxP6BLuUZZ/x/BK+7Rb7DiS53M1V1cxyqhIgA0cd+3Z3SLDtoGL6m14T4IpesZjnlEAIwjF1FG704AADQ8M4ODmc4dghvVdUFNLsntcwgiGpq5MYQkAEJDVzBEUyHdFNwREdwh2IeTaoqIgAB2pBeQuBGQsQs5lyMaOjCEBWzvpgWAwBI/1K3qzPOOOOMM74eZwL6jDPOOOPtwhHNvOnbzz7/vLJ91KZp265tU9fHugpVHHQaNOpLQcFy37lmIWdGHlgzM0IgAnfNqQNAcCA0BHSzUkrbteZbmpK7CY/VkXjLKwL46MSBh76+mbVt33S9I6WSEagKvdtR3UxEiDSYZuRhlAIA5jbUWg4Kl+FH35OZugMRmamDMbGZFs0HHQybKgKISNM0XdeafUP15e8L31ba/KYr3I7JTqnpgWYtrx/kvPpQrxFLH+2Z4dY840RreBQoHaVFeOSrzQ0BD6Ln4T33o3vGK7Tbp38ezaOPxz+S07cs9eCxMnLY/gL566ClmHsxL2qp6/rd1lRDCESDiQCHEEIVCaBtu+1ms9tuVcL0/v3ApO2+jtEAuJ5UsfK+Y5a6qgIAEVb37l10zZNmU0p2RI9VSmnwlHjtZb9tFzQZ/vZXX717ufjhBz/jvlFX8M0qTL7/8Q//+ZO03V6XriWu8qzM58vter3f7trdvqRuurznHHe7veVSmuambSeT6eXl5eX7j55d79rdRktR94cfvL/puuvnz9q2qarq/ruPilnX96q+a3vXJCLT6UU1vZTtrlj66fdWnz27/PzZ1Wb/rdMIEWAxm/7Zn3z853/y/Uf3Fhez+v5qGkP47WefG4X58mIynXS7K0u9iFSzeZwteTKfVbOy22xv1u1uO53PZotlFaq0bz/79a+a/c1kGu/ff3Bx+WC73t48e+yuFxeLWMtnn386qasYQp/61LYhhnpSi1t78+Srz36JBjK/9+mvN//pr37x+Lp5Ey6dieuqMlURRgZFCJOq7btQVVVV1yG0Keeup5K63T7WUyJaXdzLqQvMroquDpbVmrbrum65mLshABJJKaXvWhTBEEsuk0ldxZpZAMF+F63uC3fcd4Bxjs6P12ngbg5306HIIAgLIZqBGyEGYQJmxBA4MAfGwFRHrkMgMGGUwdKJQHMmZxIyc9NiJQchESIiMwdwYnbHnIqaERIxj/GDZiwyJAS4uyEyD+w0IXpKydyLFmSWqkrr7stnz3d9r2f2+Ywz7uBb3RDf8d1DRKra7Juua7uuF9Vipm74EgF9/DZ/5X4QAE5L2XDsTJh7LiUf+jkIAMeeJRqCo4Eequte3OlJqqEDGJgDuYO6gRqYFU8JQIYCDXRij8IxDBUeJIRMKEIxCA3rDBndBCxCTIjAQzkegFpR4t5kb9RLrAEznS04zjjjjDPeLs4E9BlnnHHG2wWCs6AmB1XXZNph6Vh7hsyOpA4EhDiUSquZaw4BKAqjC6EwEfFo2ydjHtRQ9siDlQZojJxy6ZNKkBgkhLHw+rQViIfKRgDEIcMcU0pt1wGSggNgKYZ+zD0/2PWaFS1EjIdd2sGRgxAlCCK6QynZHUIQ1aJaCMnhpDQSEQwIsRTtu5RzcTtcnhEvkzi/46Dr60mgfwG79HUrvMFuX+Bn3xwn/hWno8FX7QbvGGUcimnxYJUyroQnhPaBcH5ROH037ewFNeYp7/yaszky4XcYtAPMoGgppYC7CPN0SpabfVP6olpMS9/3AFBSZmY0E5K6qi8uLqIIARjAl4+/vP/ofWCmEEJVz2azruu6tq1yxsrraiISwRTMoE/gPnhRvwkc4Pl6/w+/efK3v7n+P350AborWrq+zTktLy737T6lZJq7Zr+6uHSH1PV92zS7EGeLUIXapqnt0MytRMGqrjLixTuP6ukk982zZ0+pmkynkwXRVnEAACAASURBVLapN33bts1mc3OxWrUp7/ZN7tuuywDAETjIpA777fX9GfzJRw8er9v//vefflt6dLmYf/yDD//9X/7k3/zw/YdzDJGylr5tqipwnMRIJXeb7UYkBuFifr2+qUohgNI2uaiEygC5rnNK66unqW9mi8X9B/frulpfXz17/oQQ7j14MJ/N+qbJ7e7RvXta8nq/S20jzPMgKXftbj2bVZXMfrm2n//q6f/89PEbaowHFxhVizEuF9ViOdvvd33OKZectRRjCgBQtKgpEKlDTqmkQsFz7kvqBwPxIGGfdl3bynQGQKqmZjFWXoqnxETr6/W91WWoKndIOeG3u8ZvhVkdbp2v5X4ckUbOBVEAhSgIEeCQNBiYg1AgCMwxiObezQDY1Yq6uUEQ9DgmlYK7IRi5opm6GTEhOqATEjNL4GHaqariULmvWszcnWKsRMjdzcogo0bmGGJS2+zbJ1frrk/+dY+KM87414Y/2K0wyguYHKDknEvJJTtCMbO7BLQD+CEIAk/6Di/tEOFupdSw8WDvBofKIzr6gqEBAL6SeoZDldixp+qO7owYRNBA0AWRAQRRCImQCZghCoXAA/ssCETAhCJAiERIMnjXASKgjx0TBzfwYlYcuuLJGYjXk+m0+c4u9RlnnHHGGa/EmYA+44wzzni7IHAyC0HuXyxDyp665WSOPgMAEgZCtSLMQcTcSykp56qOTGg5MSIzEdJgdEBE5p5zBgAiCiyqyUoKIeaiTZdpOp/NtiGEgYC+5XRHBfQggh6ZZWIqpZSSSQKxmEGf8kEaMm5LWBzA3UWIBtuHQZkHZu7mjgaAPkQLDvbEWopqAQBmIiZ3d1M3Y2RHBh8cRAEAT7Qzd2vNX7HwW+BraMZXkSCvFhe/cRteu+GrX9ByctBvhRcVxC8tP3LM7kfC2H3MAMTBr3vwaRxMGw9OG0exkcFxdPaas7o7zryjer7LNp+0EeFuVuILcCcmjtGrKvUJc0Fm05JzSTmnnOKkCiFMJnXRjESIaKamWlUVE2EpoAV8cIAxFEEJYKN7NICaGZrR0aP8zdCk8punm7/6xW8/ejj73qIiL91ue0MYp5PZbAmwsdLntM+5khhmizm5ac679c10dblaLfJkur6+NktNv+fdeh5inE0BzVxzTrv11WKxXC0XbrrbbDbrmxhD4FDFkFNHzEUz5TaK1zWXHuo+f3Rv+rMfffDVs/WXz7e5vGnpgDB9+N47//u//clf/OSjB8s4iV60v1rvUX0+nzF7addd12uxMJmQCIJbSe3VE2IEYKziNIT5xb3c9u36um22EvDiwYP5apm7dnv9fH9zff/996f3Hrjp9ubzeQhk/b7Z9V0jUdq+p2ltuW+7FgI3WP38V1/+/JMvrrf9G7bfzVNKqU8ubqpd2+63G0JmEjdXNQkSYoyC1WRCEkgk59Q1WwsyrWPXdeAwfP6DCLgTC4krQDYFQhJBRCvKwm3XeawQgYbK7DfFKx9c3wF81D4feJ8X9o4+WHAIUSCKzNEpEAYmHDzeAQmBEQgQHVw1p0TglXBRNS3g5lYhsBCSiDASIThosVLUTFlYhEWQmSVIjKGUgkjTyYSZ3SElMFMimk5rRGrb1tzMzcxCXVfV7EnbPrtZP1/vkgLCOYTwjH/l+COaf2Ecu3Omqmokbm5+1/7eHe3gmzHGTozeWndwVDafbOi30mY3xDEldnz5wAIfgQfd9OEQjojoSOAETmCBaBKDUAjogSBKiCKRSQIFocAkjCIgzEIo6KPPM/ugtGCmoRN05LyH3oCBKXhG1Lb0fVGm1dNqN919h9f5jDPOOOOMl3EmoM8444wz3i4G6XFgrqKwi6lEZiYCwoEPNrDBKDmnhEShirGqCaG4CRGLAAnA6IpA7iQBjipmJR8y/RyoBqxX9XQjEuhQSHhgMY6kIyABAKiquK9WKw6xAIhEcyhZedBVA9jgCTgkDRIyi7v1JQ17jDGYmZkxj14dA6GppgDVQeziDmaqhBRETB3Micjdc86p7+GbMtCPJhJvthqcnPKrPQtfPwR8HeuNd3+9K+c9DsrubHzLGR2JWoeDjaK/sPLLh3m5jfiK3+/EAY3/HUXOw8hveMMRBhOUYRQ45LoNptyjLPrwhx+jB8EP2ml84ezGgaI7uA1OkuO/gXiCW67ZRxvp0YXDT/cwnMd4VPDh2O5OzCEghTAMeN2cmEEEmQGglGKqw0iYiC4uLgHRS9E+9V2XUl/XdahrDKJubdepFTQzM0AMIi+WBHwt1OBq0/z8nz7/0+8/vPjTdyrBvttbSUt8uJgvhKDbr3Nq1+vrup4tl6uKeLO56dtdPZ3E2VymVd/1jfVt3+rm2kI1Xy61RJlMgKjZ7xi9mswvVhduur5+vt9tYjUBc0IMMabU5dwBlRAl1rHu9Z1F/On71ZOPP2q6T663jb6ZGfRyMfv4f/nwZ3/6g/fuz+vgjN7l3DXttJ6GECw1/e6m73OYXIR6GghBU8ltv1tn1Wq+ml48CPW0itX68ZfddouEy4vV4nKlZk27K6kVpsXFBbBst5tmv39079JK3+xuck7TxQMI7ABt1zU5hXry66+6v/rlF598/jy/MRM5xKwiYk65gaRmoFaFwDRMaxmIAGOoI4cqG7CIe8mpQRO1FYswB3QChyqEwILI6qWoF1MWYRYAcnNEGiyWmSgIv8rw9OvxXVLPhz2OTwsEOFEYvgxjgigc3AUB3E3NAFCcjdUcwMGSZmQCIuhTz4DDA5mJ3U0NyBhRYKydtxCiBA6Bx0BZQmYmIkIcKutVdbjTh9oXM2PGqgrWl+Hog8qx7XPT515BffRm9bdwoc44448b35Z3fn0P5LuDAzBzXVcSQghSV7GYmY0KaHQYfpgfeeGXNM63f7/4fFJVVR2UE7deGnZqAu/gjoSutzKJkYbGY7IFAAAScggcA4sIOrkB2NDCIRkbXN3QbdBYOwMB06B3BvAhrfDYF2Om4YkWhh44uoInxORdq66mzyefSVh+t5f6jDPOOOOMF3AmoM8444wz3i4MARiQiTlIjKZ1kMDER3LVD/IQNWJSRmSJBGasgOhIiHyg9oZAFwAAcC9qZu4O6GAO5k4GauiINoY+3RK4t1WVAA5g5gg4n81JoroDsztoMSEZ2laKalFEQCImBEA15UIDzyjCo8hlICkQWUaWcCDGzd1NzU1LIaQqRlNzc0Q0s67rcSiJfJ3W9tDsr7UiPjK8o9HE8STvelWMeFmi+/qDft2CYQne/oIHgeJoeOF4bPpx+AV4dxB3x+7irsvGS4c+ZZiPy0f++GAWi3cJ44F4hgOFNPoqDzJoJh4SJg+vHxRI4wdsSA06actd1t3HiQU31ZxzzrnkrKru4P5KcnH0i757ZsdDIxH1JXd9MnAOjMTEEkOs6moyX3CIrVrTNPv9fgVDXKFUVdWF0OSs7sWs6xMRhxCZeaju7fpOS6HhfGRgz15UkX492j7/9qvr//HLLz/+4OHqXsXQdO0e1vzo0buzanVtebvbliZFCfPFMjC1qS0llW6/3wiGyXQ2VW373lLfP3/61cVqicJhOotVtX725MmTZ/fv43y5uLx3sd9d933b9wlQQogSBZhS33RNk3qqp7PVsg69O9q/+8lHnz153qe8a9M3fo6F6AcfPPrJD97/4MEseIo4tZLBvK6ri9US3XLfeS5RQj2dz+YL0tRv97nZltTt922op7PZJC6X+y8f565D5tl0uby8IOFnT583u22cTCbz+Xyx3N7crJ88EZHlvfvr6yeas5pykPfefWd7fX119bRXzLz6r7/4h3/49NnVtntzPgYBB5akdOteS11PVsvV/vrK1dwUEEopfd9HwZyzdr2aDTXXSMgiF5eXqe8ZgQDAnJFNPfW5TxmRQowwmh2H3b75+OMfxemM8ZrfKKvypI1vTdh4fPzh6d93VnB0RzcapioBXG1wRiIEB1dTd3VwJ+AYEMlMCYlIAgcZbwofC2JwmFZyZq6qKCKDPhJgoObZ2ckNEc1crSAAETEP3wgwTBoxMyIBcTHYN/2+S9lAEew2j+CMM/748Yf6tL7SleLri7S+PRCZOIQQq6qqqphSjBW7mzkBjC4cgEOJ27jBoaf2ShH0yQoOiKpaShHmMd5wmKQyu81hdnfTnA4iicN0t+O4gvvwwx3QkYberDnQwfHDfbAHGVcaOsk4CK1xdHxGJCQfFdCIiCgig1giiggzoBu64P/L3pttSZJc12JnMDN3jzGHyqruRmEgQAAiuUheXVF61Jv0XdL36B+0pAdpaXFhXV7xiiQIECCGHmrMIQYfzOycowdzj8yqrm6iARTQEn2vGjIjIzwszCM8zfbZZ2+MAncxi/Hw4dbZi9/bPM+YMWPGjHdhJqBnzJgx4/3CzMBYjMA7pgY0Azkz0izEjMzEXNzpPNSsagZEAJoBTTRnVbRcDqRmOUtOCQBK1lMSEVUml3LuY67WfLM7DFkHgwSlSxsBoORKlT2MqIkKAjjmUAUKgZ2POYoYGHp2jhwyx2GIMU7MHeScnVHTBClegUTOOWY2MxEVySU+rjg8mFme8mdyzmbmiLlQsIaStW0HIp7omy+SJp/2XQ+pQ4R3iHFsuv1E+N73eGKRfMMUwv7G073JcX+O/S1/35YknZ5q2o2NXC7hg4NMlPD0FA9ExyeqfOpdfbC9u/dOeUBrP+CK78fMVIjkkgRZRoFURoYAJX6HsASIMZf9YHkAE9F0vxJQX6IlC6usKiaqKvpmL+39DBSSWkXZUSGv1QxVzRDsZPz91iMezq+pmZoCoQ8VO/EhpOBTl45dK8PACMwcQoAxXQ2cc977FKMM0TmWnF+/es1Nbcxhs16jte2h67p6GGpVBjo7O+tvXqskIjbR/X6fs3wlMZkadEP++5/8+i+++/Sj8299cH5x9+xfPVa5v11tzi4fX72+uXFEw3F3RKya5fnV49cvnh33u/bQolu4qtpenLPzr1+9ire7j5nOPvzG6vzSUgblF598fLe/4wCr1fKjb37z5YsX3eEYQlhvVvXZ+WF/bA93Q3sQMbNmvV6HRhLsrrr01z/49v44dMOr/KU6YiY62yz/6z//7g++ebEmqZFJsD30iyZcXmwtDXe3t0N3DKFebs41NE1VHV6+2r34pGuPCWi5OduenQVLw2e/3r2+iVGqxXJ58ag629z9+uf5eHDsF6vt5aPLw931608/SUN/dfUIq5p9E6oGOHkfdrvdi9fPDRCa8x9/Fv/3v/v5J6/2v5l0+3QKNKZ4OO6f1L5xngBzGg3wmYgRUhwkxcM+rTbnZ9tHn3z6KZo1y6X3AZxno+C8pdjv97d3u8vLq7BY0BBN5Wx71g+DKJBzMauoMhIBmKrpl3ZKvAPvRaI4XWOm1oGHl5bpWQmAQVGSJKSqQYCUkg8+BB+cR1DTlCUDYWAHAAbGiFMeFzlmJgQAdm4ioK1Ek5ZLWkq573tmQqydY2ICAMcuxphSyjmHEOq6EZGUBtHMjuq6Aeej8bHPu8Px0HYZQEZSa6agZ/x/An+AN+pXeorf23iISFUJKYSqCk0VuqZaDDF7FxwCINJkvgwAopZFpwYpKmKH04LwBDUBMCJWLbkgZGDTghPMoFjPA+Bo5kFoKpIyUgcAozzCcHSJxqJqGBlnMYtZ+5g9YE2jVkOUmMmQkZgdOUdV5arATMDFH46AmJwjJCAyRwhgRBhCQAAV9cyOQUUZgYmWi6ppe0n00Uc/2u8//H3N9owZM2bMeCdmAnrGjBkz3i9UjSQloLbrU2p16NkQFU0MiQBRwbKKqjKNNCOYAmS0JJJEspbYLC2OfGVZXzYKWJb52WIW0Wwp5RST5Gyjy/IoZ0EAeMC/jgMTOe4PSZWrKhdjZoPEgZFFNaWYcyaioouFIi3MZGiAQKqSMwComaqKyD0BDWAAJaWw9GgDgGBGMwBDoBhjzmK/aZ7aabdDACeR8cjP4KQrtnv178TTnh6PD8lfM1CcaFV2DhGLpPxE8wJisU496YunoxZNDVIxVRmHMXpcjOKbkyD8noAeRzFqjh9gOpmnb+9frd2/0Aev8/7VokEZItKJ0p4I5dNRpkdAuRfRyN0boOroz1iIYCmapZzyCBERFS3ZfQ9Ow/1zwdQDK5LNFBHKqy4NspPtyFvvOHh7L22aR0twU1NV8z4gIoAqmIgM7ZEcOeYQqvEh3meV4/G4299dLhpCLB27wzBUzmtMqe/dYoWIKmq58Nd4dratqvCVpK0AkFWfvd7/7X/52ZNNtfrBZVg0OQ93dzdDyqFZXT15Eo+t5Ny3eyRcrzdps97dSNcOmKwKgZCaZrlZx9th2N/d1duzZrV2zSJ1aXt+2Xe7u5vbnIZmtT6/uHTkJGlOeXe7UzPPAatlHLJmUsU6VOeb1XGIP3x6+fzV1bEbnt/sv+jTgwhNHf76z3/4F997+s1Hm7NVtVmtHWJwjlRTe+y7Y993zD5UC3ZeJO9vr7vDLscBTDdnF2fnF6zy+rNPDvsjclUv181ihQDdzXW72/fHzjeLsFi4qiaw2rHDikMFISRRF+pme765uvrkF/+qOWG1fN3a//H3v/jl8307/Ibpg2++HCIgYEfE1HWtqjh23jkCU0mgyi44570Ly+Xq7vaQ4rBy3vlwd32z299VROvl6my7ZaJ4OOSuJbBh6GOMilA3zebs7PLysuv6bMaAdV19dQuO94H7WNC3MH6GARCAERyhIzIVtfFqYGZqwgjEzAyufDYJihiwBNs6R8E7x85AnSPnmAnA0EwQwUxUwUwAhIiIQMslwyBpUlNmUiUAK9mz5aJjCpIlZe2Vj4PtDu2xH2QmnmfMAPg6fA6Ko1H5IuUUY1JTACi/fAFAHxDQauMqEpEQtfDLZvpmIcxUBQCYTURUlZntgYP9uJ6xUxjhqIcouoSp9P729fZ0k6oNQ+rNXM6CFhE8YYedZ/LMpY/DMwbPwROhOYKSxeocMyMxMoMfC/XofSIEMJPsPaOZICH4CtCDkTLiz364/t4/v8cTMGPGjBkzZgJ6xowZM943VFUQZYj73c7FHQx7VAIFk1EsnFRSTiLivXOOiVglI4pjFU2SU05ZsmRRKF3PRFIW/d6VB6gZqKEhmoIJmODEX5wkvp93e1DR4/HYp0QhKBQK0LyrCCmlJJJVywgLM+i5JLkhABkimqqojuE1as45IrTRCBjKtgSBRvqXQCWjKSF3/ZBSelcG+hdh1BtP3HI5KgFg0f9qEe/QyAcXw4Vp94MIwIRMTMyIVno4wUDNnPdEaGr3/O6k9ykOIfccNCIiEDOOXqhqADARzTR6C05HIJz0PKN2eORnT9QtwKiMB5g6V0fYqchwIr6nqsTEMGMxlrh3OCxTND7OTpUGfJP/HQPtR6dnK14aqiqmOecU4/gnpZhSSsnK+2168vvJGN8EE91dGnXREIEIFIohIxSbxmkAb+8wcRKym47FFSSqq6qqHDsuSWhxiCZqIiaSJeecvfPMDGCOebVcWekJSKk/HFUlRpOcEUGZuq5LKTEaERO7pmm8H9XavznUoI35x7/87NtPNt++WvxXT66036Why8fDkv3Fo0fHsNvd3sahI9Wl98tmmaJm2atojkN7ONTL1XqzlZy6oRuOu35XNcvtYrUiM5O+P94eNblQhapeb13sY8qpPd4ws3euciG4ustyPOyY0Tn+8Gzl/GJ3HO4Ow+2h61N+57Cr4D+6uvibv/z+D//k6ZPL1cITO7doguVD7g/toQcmJBeaZWiWAHC4fhn7FvJAvl7Ui/OzLYK1u91+d9dH2V5tlpstI8Z2l2O/Px6AuGoWwfs4tMfDbuhadA4JY4yHrvNVs96cmdhhv885D5p//tnN3/6Xn90e4m9oXf3m+wS994TZOVfXVYyDiDCz9x7AUowppsoHQgZAdi5nSTGlKovq0A+SM1WBCFKKYJpjH/s2xmGIg5khkgGIigteQVWteE181UG+D+CDi7Z97iOEAGiABEzoiBwRqJohYyFYVBWYiYm8I0YjMyQgAmYsgbfOkfMcnFPLhWJ2rtimlo9J6X1Hdjx5K0kZkKoWq43ivCEiiAhqKgqGKtCLdsrHQe+ObdsPeroIzpjx7w7vwUDjd8OY4KCaUx6GPqWcc1YwMTW1cmG592vDKTpivKq8o+9GVQGMmYvmgIhGAhphqnsDAIqMkYCoUGrdJ7HCl41WTZJkhGRqoIKWAQjMEThmz+SYnIPg2DsmUCZ0TFVwjhkJmZAdeTcS0OzGbrGhd44JURGRgg0sKRur5bz5n/+n3/uUz5gxY8aMNzAT0DNmzJjxnmEGCv3Q3V33HG9dPBCyZYtDGik9oqxZNOcQHDsmNM0GgigG2UzGyBYoXg05ZYt9n3NGxKaqmqby3omaZvV4XjusHXlCAlMQGF04bPJ1OO2HTM1MdeiHNAzITg00iffCzIWLQYA8ejEoEKoBIIrkInplZmbKJbzGVEQRUaXIZExViZjZ5SyI6ByrZDAj1CGmlLVsdv6tucMHf6gQzwBIzOy4cL5EBARI5L0f20VPXaM87p2ImImYxjh0RmJmZhYVRPTOjSNRKEFZCKND9xsyHrDCegNYidrCKemxeB2O4x0fV3SKaloobwBEQ0QwKKLdqd8UAMzGwEArMm8rj32jbX1S+k4R8zqOFMezOt3PpjM96s1HpXbxegUwhWkMiKCGCARAVM6V09KCL7nYcbyld8ITgEZqHApZZScbR0TDt52933GWy6lDQFADUlNFAO+9KKNzEmMpgRR7kSwiIj74EAKZIVhdN9vtthMZBdw5I6JkKea/onI8Hg1sKplgTqk8xVeFAby42f/TL559/+nF9z760+XaGVzHlFKMhLDarmPsY3sc+l3Lrjm/Wq63hjy0x2Ho460C0nKz3l5e8GGfh27/+gWIbS8/xNVKh43GY9e1x/2+WZ1VzZI4xNsbjT0xGdSurupmQbF7/Xo/dLlpmu1qXdV4/M7jZ9f7X7+4+eTVzeeLOER4vln++fe/+Vc/ePr0g8ttU5EJEBAbokgelLBpzpx5Xy3IhdS3x9vrOLTNcrXcXC5qHxzubq53u7uYpFqsV2cXVb0Yjnft/tY0R9XlerNYrxzDcNgd7u5Syou6do73+13b92ebrXfh9vpGRQGrZ9fd3//0+U9/9WJIX5l+xhKX5z1BP30UrYjsmElEhjjkLMRMRKV+Uio9ZppTNjPnXKgCMXXdUSQDcs4ppWhmTIRoKcZj2w7D4LwnZtXJcObrAQScLh8AAPdhX2gIwEiVD44ZzBCZEKE0c0w1LCL0zIxGJqeyVQiu9h5BAQSQzIpGmcyMGZumRrRC1gRzVRVkbIjombmkihFySSaE6VMc87Df76uqclVF6NVgiHl37I59jwBgD4WVM2b8u8LX6HpyAhGbWRxi17bH9ui8l7Jmg7G7AsYC931Nviig33UwMzMVIeZSm9fpSl8cwIoNtGQtiwTnGCZN9OeBb1LchBjYV8wVE6M6NIfGOBLNjpAZmTAEX1eBwAiN8ORKxmCggskMUIvDPQIgAYEiGpbLaBgSB3EuUe39b5yQO2PGjBkzflvMBPSMGTNmvF8gIZtS8JtV44aM3pjIBHKdCYspLxqaISBN1CkImCgIgCBYcfgFQNXS5iiyXJRQF+/YO2bCLEosoVg432s9T36mby/2JUvmZGbE5IkUydSK099J9Fv4RSJGI1UzEyIqdAQAlCyY4uZragqKCDmLmY7hhKAKoiIAAGolFlEBSnQifAVKYjJEnaTIJ3H3vT6YyE5GHDhqbyb5zrgLEtMSqYhUtDFECGYmZqOH8xhWU2yj8SEXZWAASFT2TnZPsRoYgGqJ5TulD44CYwUtQfL3r+NEVE+EUAn/O9G3EzE9cU2jmPleu1uy/swM1MDwgd3Fva66qJwmCTUUA5DTeCdWupRGTEGLWQqzK29XFTHRjHksJ6iOr3oCTVN0v1XFB5Ybpyn4YuPX6VwWWh7AQEWSSN/r5tGjrCIiIVTMjMzAXFXV1aMrdgwpFRY95xx8YEDv/XKzefnZp1VV+bpGRBsGybmuazaTnCXG19ev+2HQ34oLiNl++fz2737yyQ++/fg//ukHDaHd3Qx9+/L5px989I3lcjns913XHXY7qFfNauu27lZyP/Sxb/c7JkfLzbpe1C8/+7Q9HIiDq5arxfL88lKlP7TH/eEA5HntC6u/WDYEI5/onNuEZc7peOxAIcfBsz1e8Q++cfmr5x++utlFUX1zH18H9/SDy7/5y+9/+8PzZeUcoyNXeby9edHtb1G1rhbkggOPxEPfd7s9AjSL5dnFo+3ZBVu+ff7r/e11P6Sw3Dz56Jvrqyfd/q477lPsiXGx2Sw3Z1VTo8nQHkR0e35xdnlBlX/x6acCTC70cbi9eX22Pb/u7Wf/9PMf/eOv9t27tHNfChvfJUiEaBBjbztp9wcEKBmnhRh1zi2axnl37Noh9lUVyAIBgRkROe9DVdVNXVVVlkRsiMZMdeXZkapIjjmltm1DqAwwpVSaS/7o+MILN97/TwBM7Ng5RFAzsOILP5VdSklrvBQ5x8Fz5dkxESMBMCM7YnPE5DybZjN0rgJQ0Swxl0Jd+SAz8+mXSs5ZVbNkx44rlpxVNHiPiDnlXnICr0h9kpSEvvAaMGPGjD8GDEp1NoTAjgnHcnLJnzilhZqBmj2QAExLlLeAY3IxEyER6FQHO/36n6rZ8KCY/1bjVxnVwxVhWeAxUeVd5X3t2ZGd/jCZK2ICQmb0np3DUPoHCUCBkIhdcUwrycRQUjGYmLH0CBKRAoJf7GIycmEF3bF+D9M9Y8aMGTPewExAz5gxY8b7BRIp0aZpPvjg0sVKuppGnSgxj5lzyIyORbKpQgkhBFVNo7PBZMEQU8o5iYhjT0QlNK746KacfBaqanaOHJ/Eue/c/ZtBlsyJiaiua67qKJKzqCvmfeS9R9+h+wAAIABJREFUK0JbN0YHQkwJwJhJhcB4ctVDJFIQAWRkACAwBUNEV8TGAI6o7E9OHsRFyfwVBHEn74eTwNjMsgCzoREoIpNa1oSMSPdAHdlnRCyibMfkPTtyNMbwkZlJFiJix0xMTFRkzicZ8onXLRYcgMX72MzwQT6hqJZ4H3jgcKGmb0h9TgT02NN68sSA6RXeRyze888nC5B7dnrkjUFHemlsejUDA4WRL54eWqoIhDDJsu+PbtM+0BCQiRA9EpkomqVExRS62HybGqAVZh/AxmOOAmh409H7Ief0zgbk0XhaszKzY091LUPXtV2MajEuq0rOzw5tq2Cpa0mEEF+/vl4CbVZrzHLY7/t+CEhWaiHO1fVif3u3XHfrc2AfHj169PqTrt3vrYq1r5Ccc/63c1dQgNe74z/+6sWP/uX5xfn2W5dnTda7V8/a3e6uqpbLzeMPProN9e5mv7u5iX1crFaPHl9lU2r7PAyH27u6DovVcrM93+/37bFzfMNmy9WiObus22O7v03p0LfG5JfLsFif9/2wvz3c7m6P7fHs0cV6vWkW66HvD7triQfM+PQ8/IcffvsXn7785NXN8MCIgxAfX55//zvf+M6HF5uKF4GWlQONx93L6+fPEF1dr8EtBX1VUe7bbn/XtQfy9dWTq9V2C5p3r153hztEWK7Xy4sn68srOe4P1y+7w05F0FcfPf1WVdfxuLt5+ez21avt2UWzXAnQ9fXNsxcvvvfd7/uqGo77KlRGzY8/fv63//z8p5/c/Pa6MoT22J6tyLNHRGQytTREE60WixBCXddd193d3dXnl4vFIh76KGqYCdQRioioElGofM65cr50iCPhdntmBof9fhj6qq5TisQeAXNKXxMN9DtHUSpOJQKAERnQEXtmGaIZcEDniJkIjaBQPwKoZOpcqEOogmMCAGVm58j7ohdk77nvoogR1aKWcx76wTvf1LUqEFHwQYtjvEFKKcYhZ6mqyns/xMHUmrpJOXUxHvocw1IpJIEsYyfNzEHPmPH1gZk65xbLZV03oR9KSblcXHBSQIuaqL6pgD790n+IMay43NGm6OJRGV36H8AmnQBz6VApFUl7Y9GA9nDZM17igvOVD1Vw3oFn8AyelNGYjEdOGRmBGavKB8eOSEUQkZ0ncszsHBIBEYYqBO99YDAhROc4K4qvq337uus+vt5chPiHmf8ZM2bM+PeMmYCeMWPGjPcLJERgDsyLxvkEmFCNkNh5UDVTMAUmI4zZihuDqQIoABcetDicAoAxA3ojQR+IWVUKzYxoTrITxeqiWne+WRLfjuK30Sj4fqFvZiKZmZer5ePHT0om+pBSTqKijFwsVnNOKWcEcM5779q2U1XvvaqWuELnHBG3bSsihYo2syy5bDqQgImIOKWEQD4EkSyaJUsbBkaKQyvyZTmEOI56VORYMRoGtNJJSQQiYKpEpKaEQIB6r4meHKHx4QHFcc5UFLuFpAaDlHMpBej9TokmJfSJocbS6T+OxCYR72kPhYinpMEx6w9sJKBH6nliYkZq2x7s1B7cYfpbXvVEQeM9QU3TkaejTKpoUDAzw3vP1dGQA0GLAcUDKujErI+TAyMjrmZE5J0HA1AwVROFU2BiOV6Rl0/ZjipaJlSKw8e9fvudGF1HtMi0kUw1DoOKVFWllpGo67vd7m5I2Qw4BNOiuJTydM67uq6rqlIAYFaz3HbMvD07q5cLYDbCIcZhGADAO0cAq+W6JGR+8ai+DEPSz14ffvSPv/zu08fbxePLZrU5O797/XJ3exeHvFiuzq8eZ8WbV9dd16vpebi8vLjc+/1+f8yx393cmEqzWBjS3e3u7vZ1zinmbdXUTz765vULjH2bY09ekT0isvccPHRDP8T2eFwsl45dYlYAUw1MFwv33Sfb//avftD96B9e3uzyJC/erBbf/daHf/Gn3/6Tjx4/udjUjNIfuuPueHjtiYB806zW621MQ3c8SN+ZSt00dbNomkV/OOxvX++vX+Ruf35xWa3OOFSHu1uNvcQeEKvF6vzqERL0Q9u2+7brQl1vLi6zaNd3hnT14Uebs3PIucvWd/HjXf9//v3P//EXL47xt+SfEbGcNe8cQlK19WrV7/aIlHOGlKqqPh6PKtUZYqjreDx0faciPlSOCMB8cKJybI8imlJ03rPjuq6G4WgmVeUzIiDEYcg5B/Yn056vEx42syhPgkRPVDEFZkfkiH0IDMA0fjC9c1hyBhSQwBE6Lm0QI1lUKoCqOaXsHDM3AKaq5VMDRjDa7JBzwUz7fiiXx/L8zgWzlLMej23fdZJyCS7MBpH8UYbrFHdD7gSSgcIUNjZjxow/OhCY2HtfCnhNUyNRWU+UtUP59yEBDQBmbHafR/EAWpYfbxLQ995dUy2cRxN5ExNBgxzfUCGYvWPRgIjMXEpqhURmQuc4MDgE73Bs+AMjtMqTZ2Ay9MVyTJjRMTiHWBq/UhQlEucZHTMDmRiCVQ480fcBWp4tOGbMmDHjvWMmoGfMmDHjPcOIUIAC+YDgkR0SICGxMy2UoRiCgikWO14CQzO0or81Ezk5NDggQiMFBkMFLqo0ZjRygEY+sA/guGTgjRTlpKrF0XdhNGh23o9GEGaFOFURdsQEhACmJhmJwASMygDBtKieJQsA0NhfbaXV0QxIEZAAzEAQgRlVCBEdT4YQoz571PP+G6TEQ+Z85HnL3oagbHEUDBRgTBGEIrqeujtpEg/D6eUXwrT0g5oS8sTsjlLiQtAgGI4nonCyijCabzzgbyadMwAAECAUJ+iiJUI0A0MqwuE3ggTv9dCg71AL28Od23R4G21fx7Z6mNw3Tg/EsSff7ptkp2l4YJNxYp8n4bMZ4PguG509RjU0O1MzVhWnZKYjr33qwz0Jo0beHQBVafS5xi8uLNj9/5PcKcWUSxZSzjBNo5mVWyqAnHNKadE03nsyI4QS12nsiAhUQVVEgvdMXLjtGCMhcQjOO1D1PgDgOzOUfhOowe44/PMvnv34F599uA3N40VdL1eb3LXtMNyq2tnFo/XZtuv6vu2Px0OoqqpZLJcrU9jvd8fbGzIBRB/CerOJx+G422eR7fl2tVleffD05fNPJcYUE6J0zIZUhUDb7dANeUgDdeQCE2622xQ4ZjHhD4H/6rsf/euvn7X9sDt2gMhMjy+233v6+Aff+uDp48sAIN1xaA9xaIn8Zntm4OuqJpN03PXtMYtWVb1aL4OjoT0edzeHu5sUB1c19WrbrDZR9PrFMzTJObtQV6stV/XheJNil4ZIVdNUjQ/heHPTtq1frz64+qBZr9rr6z7Gm2P8u58+/7//5dPPrvfyWzGP0/UCqxBwdPJB7zwClETK4g0BCFVVVXUFACkVl3kkRMliZiraay855Ryd25TaGDOJ5MNxv9KrEJz3LucsImY6ppp+DSjoUw/7g/9P4aJgAEzoiVBLn7w6IkbgcsGz8dKHCEzoHQUu/Q1mk/d+uXSLqKqKYM65FLJSyjhZHJVvVa3cKZeQscmqKGdR1RRRkqiIZrHS1k6cRQ9d7pJGLZfmwnz/MeZxxowZ78IUPzHWwE9LpdOKaVw6TlDFkw3X24eCsthBLCnPpmZ0suswM4Bi8IVmmsXUjNk+vwB8Qw4NUwUcVCQnIDMzAWMkIzZEAkaycc1TGtYEgBCQEQBRwQCygQIwETICgjEqgTCyI2M0IFAGFgSG6psv8vPl+5zyGTNmzJgBMBPQM2bMmPHeoaboTKzQymLqkQnQckZmZFZBNTHQosn13puqisoEMymkHzMDIAKnVITGOMR+iD07V2QilcuiooXYnghogLIuP8FUjYkA4Ob6psvJVRUQpZiO+2MVQvDBe9f3fYyRnWMa6QYzIyJmZwbDMDjnvPd935uZc260uRABBAOVnJx3wXsRAwBmMhMDI+ShH2JMowv0V2MlToTsm7eCniS5fPLfQCxJg0iECIWN8t4574p9NhKGUNFEpuNJIVy4UULHDhDMQFXKMU1HfU8hunVU8U4iZZo8pwsLNBK6Bg/ck9HwAflrNN5heh33m7ZJI/zQ43dUTWv5kugUMn9v3FFw4tPNTlu5E1U+zqFNP550zyqiZS/KY7gjMzvHY+Bh0T+Pr/KkioJxyEUbPimyCwcNAIXwfejr+I5TWtIpVTWmCBgAMVShrpshi6pqSmkYRHJVVWViVTXnnLN4HwrrzcHHlExVUgIRJB5ZcSmCLEgxmtpvLW41gJjlxfXh//nJr759udiEq8eb8OjDp88//vVhv9vvdki83m4vri7vbu/6btjd7eqU19uzxXKR07C/bdvdThCWZ+er9YabzbNnz+LxuAdlwu2jy35Ix9ub3B5BB5GMzteLTb3ZVmHY314PXcc+h6Y5254NTXNsO4oZHXw70/e/8fj17b7rBwXYrpbfeXr1/W89+daT800Tht1NPt7l2BPxYvuoqhc5q5n0x1083JgI+UVYrpvVOh6ub15+1h12aLpYLlab82q5YecsHg+7W0LwVVMtVlWzPLbt/u51ip2vFquzq8Y3qT+2u11UXTTL7dVjTX3Xd7eH9pPb/kc//vUvXty1Q/635/cL5hwAzCwErxpR1YeAhKqaUsw5B7OUYl03i+XCe6+STdWRU2IzExFCTCkRKDrt+y4Ez84PMY5Xzn5IMXHlmImIypUW1OjevOiPiTcJ6LeBACeePWMSp8RETEhcLIJUgNkcYxVC5Tg4cmSoasVFBxwjgYGoMjskjCmiAQKKnAzfSUTb1OeczYyQYoxZcnEpAoSUEpgxUnDO+QoKv0ScfH3TaZ+GaCBjigD+LuWfGTNm/D5hICopxaEfhr7v+x6Z2DkiwgdGzA/TK+BB68Tn12BlCYFGMAWgmt1nEZevS7hIackaPcXgHXXqhypoA8iqfRqCZEBgFEZzBFK55NkRBE/ekXfoGIMjUwJjZAaHpVEsjdnYwOzZO1cE1EyByXHxkWMJDebBgD77yTpefi0u/jNmzJjx/2/MBPSMGTNmvF9IFkTd3XW//tWvoH2d9y9BjQAdkZoCgvM+5jjEwUyZyDsnIqMZNI/sac45p1y8FEr8GjGJSc4xSyzsK7NrtsfXz69Te4ScP0dejNJUVRPJJWuLmHTQruvIeRE1wJiyqmVREVVDNNDCA5ohICpkSQCIxCnLEFPhKkurJgDoGC7H7JGIDVhN1FRUSuy4gmUxkRJvQwBfHvk1qWRBi7D6gafwSRpcqM+RRh3547L/kSwqRIQjHaxlJCVVr3AoiGgyRSKeAASAAw7MjghFZSJeiwkzkmHpiDe91yOjYpEJ3xPMk6D4/sD3CuDTz8tYJoJ6+jEAEoIxP1RMnyh7g5Nn4z1NddoYFl783knxJJt+cO9Jjl2efhRwA+iogTJjYnDjwIgIM57iJR8SY6ZT2uEkWp0Ob1Yk2fdn6t7g0SYlPpg5pgzmHG+qbT8oquaUAayuq6qqTI2ZnfO7u9ul85V3mq3rumEYoujqkQA7cB6JUkw5ZyAC77z3+8MhDwPUqwbhcDwYaKnffNWixzSl0Cf5zz/+5Z8+ffLB+Xpduc23H8W2zzm37fHm9jUyLDcbF/j2end3vUtZiN1ytTw/v9Asu8M+H1ojZuCrs6un3/jGs2efdYeWiA39dn3O2fYxS7I8JMqWeSDyzOSci7G3nChzyuwcN1VdB1saDNp+/+nls1ev98djF/N3nj7+6z/7zl/98DsfXq6H/a0M/dB3KrlZNOvVNmXtukPOgzNBs2axWF5cLdZnKun61cvrVy/i0C6Xy4vN44vHT0RySklyCs4B8+MnHy63Z1Hk9m4fu9Ygh1AtVxsQvLl71g6DX6/W5+e0Wtz9yy+vX7347ObwDx/f/qeffnpz6H8X0tGmsoRgDo7qpvLOFXeNLKkfupQjE8UhDf2wXG6cczFnTZl8CM5FYu+cY2S0w2EnIuuzRZKsqsvVcrFYOPYpaxyS817VUsop59/u7fGHAU39EwTgmasQqhA8EQKoqJgRABMiI6E5Qu/IMxOCSoaSx0UUnAvemUHOambOoYlmyWTAxKEKcYgppRACAqhkVQUEoFKkMskJyudX1XsXQiDAkvlKTEZsHJCSAhZvIQNQVfkyT54ZM2b8QVEyhFU1phRjIs9Ztaw/cFxRQRbNYkRjlVtVzew+zvgepU6uRIRIJTDCTE/Lk6lTZex6UxVTNdUsb6/9bCK/T1VzUW37DpGEIDB4QiWwnHseSWfvyDtyDr0j58gTeRqr8mJAjOTI80AIiEU/gYzgmBwROQYOUPe7wXq0f7h6+rT6l/c46TNmzJgxAwBmAnrGjBkz3jdUBExjHm5fJWiv9XirIgjgiFUFCaq6iSn2QwdoTOSYU0yq6pB88N45MEspDkMEsJI3WNcNO86aRaNKUlADQHRJq+54AM04uXjqpIPGewcOy1liTEWJPAxDMiMvqpByRoOE2TkdtxFmqlrkz4ijMwMAOOdSSinlEAISghXlIKopFaaWoLRbiuRyKC4ErGGKJdnuywygH+B0J73X+eJJWjv6WIxmGIXRBEMyMoTSbl560c2smDnEMUhn8k8GQrp30iBi4pFMV3PeEZKalh8RU4kZnPS/k5r4vnEVR/5bYYz4Q4CixsUHCYOTSYWNcfEnnvdLJI9go6546scffZnvqeUyjpNzy8m35XR3OD1y+gqmjeU41MlBozyQiJDdqOKGsrPUafwn2+iR1LWH1B2W3eQ7T/CD2w1Mckop5wQAzBzzYGAln9ARI6FbrZxDaQ+GsFqtfN+j6nK17roeiB1gPLbd3W7ZrLBR51hSBm9q2jRNRipWj5vVuq6q31Hcqgav9uk//eTTx9vl41X45c9+hqCrzcYHbtt93+1jOq43Z2eXm5glDem436FBs1xtH38DqluVlA/dzbHnpNvzR5eXj17f3Ox2BzWAtNEk3tdYbCpB+/aQcgyhubi8PLTHw3F/2O369hiYzMwvlovV2dN68R+SIqTt0j273f93/82f/Q///X/8kw/ONB33ux2KIrrFerVcrdFy7PcmrUmOCsrV2cXjuqlid7u/fpXanXfo/Hp5dlZvt6I5xd7UEJlDc371Qb1a5ZSGdoexi4OuNmfr5TkDXl+/7sWWl483V5f1ou6fffLsX3/62cvdTz/e/W//+ecv9in9zppXImyquglWO2Pi/d2+7/vFcrXdbsJy8/Lly6zivKvqmtlV3vdEWlS3CCbJedYc267tumG/PyxWK1PNOd/e3DTLbUpCoaqqhYqcX547F8Jnd/nrykGflIkAQACO2DvvnWMALI7wUwmNcXRK9cxMiKCmgjh6qTIzIomIjrGlqCpDjGjgnSPyMUqMqbR5mCoRIuDEGt0bEJX0QmIu5UTHjoiMGJHUIJWGFwADnLo4Zg56xow/PkpzWIljVVURAQJQBRxjAMsCIIslEZqiHlS09MB97nNcCoXKREio43dv9BuNJh9UVoBqqqB2Wvy8ObhxLXGqqquZgGYFh2hlAamqClpiVgHUQAyzmhfIZGnKuFYkdsRqwiU9VUtwNiEwwdgiF4A07pJK5f/ir/6Xu7un72XGZ8yYMWPGA8wE9IwZM2a8X5ipKYiZY/Z1TbQ+uTszkXMuVJWZqo5GEIzQ971kYWbvnXeOEFU054xUKGhBYkQQE5GYZIgpJkmiVi/qRSOLZhHcjmnUnijgiQAY1+uih0MrotevXx2HCOyBo6jllNCQyTmXVUVEnePixiuiRDiGEIoCjNuSmHLhJ0+sbomLwcldWlXNoAi5wUwVcracRUUmNvM3nchxOhFK4KCN/s1kxXFCBRBBIY9iYXST9hkmakZzVslVUxfPkJgiGFQhICKopZyZGd1oYlysG6DQ94VuMQcnxvaehgaASRaMIxU+SqVH+TGKjN9NDh0EJ6J42u/B+MCR133w/hll4IhvaI8f3OetjVwZCBg8uLvZacwjbW2nmx8exyY6X200HNGp9sCIqA8sRPSUWW/FqGS69zQKnGSPb+wo75/M1CSnxDFKkpSGYYhmBAAleq4fooqCSo4x5xxCVcoaSMCOiUgKS+qcd/4uRkdQ7GfKFpqROFRVXQNzVVfF0ft3yUIzgCT2s4+f/8PV6k+/cXaxXA3H3flmtd5s2MHQt92QkWizPv/gwyevnr/q226328Vsi/X2fHsR++Nxvxv67vrVK2Rebc8euUd0fdO2bSAKIdRNQ00TQn1sd1mSDj2YrVbL1bJhhq6lnAbJ0Qyka6MB+fBkQ3/5nbOr82ag8L3vfufDs9rrILFPKS6qpq7qUAU1ub5+meKgAN6HUC+cr4m43e/aw91xdxNTXK7Xi82mXq3Y8dB3x/0+Z3Gu3l5cLpbLvu/aw21sd4h2dn65Wm9N4ObF893dgUO9vPpgdbnV2P/65z+7ud198mr/T796/c+/etVlfSfD8BtiLJepmankHHMyNec4+OCcK+/GFNN4BVDNMQ5db6qePQP1x1ayeGajoJKrqgkhmFnfd213VLO6bpyrgByzZ+ckJRVNOU1P/rWFIQADeCJPXC60aMXr2TVVBaZM5p0Pjr0jAzFTQnTO+eAZwcxKgbNcwERizhJjRIPMuXyQVaHrWkJ07KpQIUCWqCIAEELw3jvnsmQziymr5CIwRDRDTJqHnPqUkqmWItaUmDpjxow/PN7yzUDE4L33rtjpUDG+H382/osGRMDAo9MXguA7PaBLnwOSUlEejFIF/DwBDTgWgBGIwCxJevcC8L5RCpjdcrlYItRgAcEjOEQiZEbH6B17R56R0AjAe/ZModilMTvnkIgcOkfMxDyuiwiBR6KdKNTUrPv9sUcEgO3249/XnM+YMWPGjC/CTEDPmDFjxvsFIZnXxteXj66CNhgbtFEdWjS1o4hMpETzEUIToyp4H0r6NwIU7RkyAajmBKMBsRiaIQiqiKiqW17dpNfrzdaH63vngxObAwCAapCimEHw1XZ75oeUkcixqeWUR40IYvGpYMdmJlnUDBGdc5M1tTE751hUVbVwQ1AehVDkxcWaOKUMYERU7IwRMEZBi0P/JQpZgFGe+6bbw8Rj3hOaWIS2xbGCTlF/xR2ZSu5esa4mImZ1rOpCGDksZjaD4D0iApgXJSLHXNTCZvfto2X/xkgGcOLziSbl9SgFtiIqLIR1oeMfngKYGPOx0/XBqzrFAj68bfrK3nE7TLxvGR7gJFsejTcmlvh03zeI5vHrkyT69K+VLljD8f4GAMSMRBMZqKIyjmksaOjpWG8Jst88p/b29wbF24WJAaHEoFWLDRGpaoqx6zsRsZwti5oRYdd1vFp6pJwlpSQGqsreh6YhomHompWi90X6LTnjVCQQLZYyv6si1wBe37U//uWLP/nw4huP1pwhJamDr5plTFn71B+7wPV605ydn+3ZtYe+PRwQ4Gy79U3DCEemw7G7ub5m5+rF8ny7JgQ1TWkgH1yoVttKwNrumPPQd213vKvrahE40HKIPosYQFLIMWpOS5aPtv6jx+frq2/Ui0Vs72JURm5W6/Vq7cBUUt933fGIRK5q6sV6sVww4WF30+7u+vaQcw7NYvvosmpqBMj9QCrHwwHI18tmtd04tt3tbn93LTFuz7ebiytAOtze3b2+FqD15Wax2ojA7atXu/3htoOffXb4x1++vD70v7vlb3mHHI/tpskIGYDqunLem+owDBmdmUnO5Z3DzoHZ0PWsuXLOVEupjBlDCFUVmDnnnHISkb7vx6sZMQB674dhMECR/DXxgJ5ImPtrw+nG8gUBOANUQwJmYhpVjYRIoKqSk4IhoyETsys1PzDDKXd0EjKPda9yqYxxKKWuUqKj4jaEhaupSg2MiMoHHRGJGdGYwFdBTIY8HDV3KSUZC4yKOFrxfDUC+nTvr3MxYMaMrzvw5Lg8VaDZubppnHPEzEwlKGPsnZp+RZbCkcPJ7AuRaXSF/pwHtJVlA5Q81PLoqdYOAKqmp9UFIhYZhem7P9o2Nk+hgUMMhIGpZl4gBTRP6BnZ0UhAM3om53A0dyYq/zpGIiKEInlmB0RaFl7ESISOkAiNCB1BoCpw1i/3gpsxY8aMGb83zAT0jBkzZrxfsEO2KjRw/ui80sp6P3kJw0TEmSbRnJlHIYqvFBGdD1i4T1VTU1NwDKCQU9G1mQmyI+/BM4CZKlZnq2tplssSFXgybMDRXQ9Lu3ZKSshNvTg/v6yGGNXYOzCQnMvYVA0RCImYzMBUJg0xiqqI5CzOee9cFlFVMGCmKdFu9FtmJnbU94OZOcciYgpE1HXRDI7HLyJ63tyWGMDbipt7p0CbmHWE4pFBSMgwRhHCZDvBzCVrDIIDAKKST+jYOTDgqcn0ZD84KZNx5P0RS+85MU2866iJLrePguGSEz+qoXHS/05sL55IGD0Jpu9fLE6uFg+k029PypvzMBHO9zOEk9/Gg0e/pad+wGc92EU+pIdtTA4czUOQkKctbOmtFZXSjWtYMhLHWbKTAfdEg9s7Dv/GqTUDRPTe94AAEEKogkdEEUk5q+g4k4SImEWOx2P96JIB0zD0fed8BUVbXlWhCt3xYMTsvZgRooiYSk7JRHNMOeeHgY6/NZLYr57d/F//8IvvfvPxn10tU9bDsePgqnrN5nKKx90+J724fOx8TXS3v931u5sOdXW2XW+WrnLZtGsPr1/Y9uxsuV5fPrrY73Z926ZhyLU063W9XAuiHFVie9xdawxV1fiwqDZbQTKkFFN3PMbhGFiBpVm4x2eLQe3FYa+IzdnF5vwieN/vrrvjLvaRiKtmFZp11TSIOhxu2tuXQ9uBQd00i7Oz5XaVuq7bH0B10dSI2Kw26/MLZNJ8zOkgeUD2zfoiVM1ud7fb71LK67PLs4tHoHD98tWrly+pWr443v7Tx3c/+/Qm6+9B8GpgKeW73e5xCOTJTHPOYDbE2LZtQHbeDcOQciIiH0IIYRgGi31dhW1VHfsupuSnj6EsQqA7AAAgAElEQVSI5JQR0LE7Ho993+cs6EdSJucESA9SRf+YePN691A8fK9TZAMGICxVTGRCQhq7JRBVUy4f0dE3iGOMmkVNCZBxDBcAKBzNyNQg2BS4ynVdIYKIAiogsXPOOyJUVRUTVQMgJu+9ZCM08hRj7nPshPqUh8m2ye6vWr/5tNqbX//WHPTv8tg/CL7o0jhjxu8PDxXQiEjEPnhEQgDHLjhHzKUrqixhytqGDFXH8nJZl5KBqL79ltVSVp90AQiAaAZM45JKULE4ko1J2qg6Niq9c7AAYyHcITpCAvDEFXNF4AmdoxBKcqoFh57IMQbvvCMEIAJXmGgEMGVCJiBGRAPQooNmRueQiYAIHFvgJnAfbWagZ8yYMeMPg5mAnjFjxoz3C0ZUl8VILYkMJpGdRyARGY15yVREJZOxFgcGzVkkdm3ZOeQkwzAMQ4SiPDNhh0QACFlBFNCRgooZ1YdXr25TSmJmCISjGMXUJlkJAJSsGFAb9xfFFEJHk997vwUA0JK/x8xMMBk5GGIIo78oGzCzc05EwKBYBJqZivjgQyjiYqjrJuckImAkgs4Nk0/HV5zNYqR8z9KOhq9INOn/kLEE54yR7jBS6ppzdo6dZwBIMfcy+OAds5mJZDMo+u4UMxA6Zu+9iJoqlb0UkqoU40J2DgHVtIiDzJDRillqGVmRJU/uGYaTI8lDhniMAYTTa7l/jTjNzOfURvea5tG4Y5rCN487GTkDTiWBf2uibZJ9m56SFMEmOnpUSo7idiiMO6gAjMaw+s7nOMmw3/UqcDTV7rqubY9gVtXV6+ub5WrtnVuvV9WiaZoFVSEeZIgDEbF3hFh02CK6XFWOEFSz2fXNTe1DYAdZkDGEKoTKJDMR5tQ0jRt17r8rDOCuHX78yxf/649+8s3/8W/WQff7OzF5+vSj86sPX7149vLF8/7YD0N6/MHTs/Oz/5e9N9mSHEmyxWRQVQA2+BBTRha7T9fr5uHQ5OGCXHLNn+DXcMNf4Z9wxcfmO/1OVw9Z1TXlFJO7uU2ADiLChQJm5jFkeGZFdGWTdjPT0x0GKBQKM5jqlStX0GR3e7Pb3UUZ5hcXs/ni2bNn33377eruJuWhSA7domtCyWm73e37gfb7y8vLbjZ3jlLPcX+3Wa/3tJ/N85PnC25nxcwxkxbIezRF1X5z990ffxe6BYl4HxrGxtN2e3fz6kXuB++bdrFcXFyFtssp3t68urv5Lg87h355cfno2ZP51eV2t96u71If29Bstvsvnv+iWVwU0NvVDco+5+ibpptfXz17vr19c3dzu9vtm9D+xS9/Sd38m+++ff3qBSFjM//1i3/56pu7m3X8JKyaiMY4DDEiNewwl9Lf7WOKQIBoTRNiTKIaQiDE9WoFavN2FrWoAjN77xFBRFRKzhnGDxY5x7OuU9XNZh06C873fZ/zwnmvpimlPzsp+EHeFA0MCIABmNCxaxofCNnMMSFojInJvMO2cY6rw0bJuSCAllITNLi62AOQ0cFDyMyI0DnHTPX3ELyZqgkAIIP3vqYQhNCUUiwX5z0TMUHJGktKkpJINmIfiubNfp9FaljODk+Nj2J8JP4pTjlvN/ezxpl9PuMzoxZ6sENsGBFMd7sdIsWUurbNi4Voza6DwwywZjmoHGQMeAilHwocTydQNKsULxw8xKYTA8B40lppwwxApZSEIAnf5XxrlYupCTRDVRCRAkCKRqigxHXWZyJEYPUhTziWUobqv8HkmYJn79gHV5O4ao4IExAZIRgQNS10F1u1nez6z3gTzjjjjDPOOOJMQJ9xxhlnfF4YFKdsNuw3q5zXtr/rgc1A5UDnAoiimuOx/F3RJJK1lEp9lmIxphgj0WhdMO6IWNSKGiAJqJjyDGO/N5WD6/NYGe+ogKnrkOqfDFXNLEZiWVUlZwSrZ6kLiVJKlcwwM2JN7RZVQyJTrWJVAFTRXAqYjTWxzERFVFUkpYyIiCnnpCKIXIpMftf4IxfgJ/reyeTjOM5m1dgU0AxRVXmqegOjKnt0BTEAUxVRzGhqTFUtC5N0WxBJFXMpKlLvUfUVrGYjAEhqoy/HqA6Gg7/GZHdyIIZHGXrtwlHGjPc4aJykyiNjPlHZR5uNo/ZxvHqctNhHAvog4saDATOOymQ72JZMortT/nu0vDYzA0WbappNNtUGU83Dar+ikyS/EsHjuNUhVjv4TU/vtw/DLJfCJsF7UzTRxnl2vhQZhni7WV+t75Zt45qGiO9Wqy8uHzExoTVdu1wuDUC9VyLb7Np2ZjkN+z4M0V02McZqFgBmkmV1t+77QeRPdoUAAABRWO3S3/3j7/+7v3r+v/xPf/30aXf35tX6zXo5m88ulos47NbrYbtZ395cXF4/evLYe7pb3eb9DsE8UbNYPnr2xN2t4zC8ef2qbTdXjx4tl3P2/nZ1V0oahv1s1rZt4x16H/p+JyX3Kb169b0CIjEC1WTpmHLKmTyy5BKHq8urJni0sn7x+812W7I2y8vZ8pFr5t3ja+o3d6+/efHtH4oJEHZXi9nlJTPdvfym3+/ZcDFfhm4R2i50TZG0vrt59fKFI1jMl08eP/bd/M2r7/eruzQMF5fXj5//gmaz7777/c3rFyYKYfbVH27+/qtvvn2zKZ+OVkPk+XymKjGKqqlo6uNiNm+bBgBSGuoDJ+ccQUpKBuqc894BADOmlLzn0DREHELoZrMhDqrWNC0RhRBC0+Q0NN73ux37EFPKJX+KOMXnQn26MCCP7sqjU5Gq2GRHpAqqUGocsGShMY2mPtWZakoBuZoXwgagqoKEzBgaX8vGihRk9MFX1v7gtTMqxomcd4QGJmY1HYdCaJswk9kF3eX1dldEal4O4I9yNTmTsmec8QlxL56FiGYwxFhyub292e/2MSY1Q0cAOFZxRqzJXvcJ6CPvfBoeQlMYCyRXY5+JQNbxWKoPEJtIcDSps853SwTY8Uz1hxpk0YToABSQCZyiAPiCTOaZPKMjLN4FD0jmiDJLZg6Og/NFwLG5IoiAaMxMTIRAqAhmgNwKFd73MSkAwD/8w+e6B2ecccYZZxxwJqDPOOOMMz4vyKxoNMnb1S3v3+j2TYoiYohcVaxoSoAO0bNHQgMQTapZNTvvmB0ASxYrhZzDqvgspmhqpogGqNXl1oTcAiSTHawpAI6U82EBYQCGBFUfJ6VkQ9FRhc2ERFhKqVmMw5AAgJmZCBArBWmqSKPcWEQqEVtyqXtW1bZoIURmFlVEZB5SimbiOOSkORdT+CkKNUQkhGp8gWN19Uoqi4zJoVYlfoieGQG1VqUbfYFHl0PE8TJFxBEdZMJEVAvcGUDOebIuNERQhUqzIkCZvGKPfPGkVj5y4pOpx8QS2wmLjKc7II6uy4cjJkfW+vvh58G4Y1RWT2eyw+84XjsA4XHlWHnydxXTeNLgVJTeCECgLh5V1URtsnCsfLNIUVFRtepDrmaqdmjiwHYfL/fARx9vNzM5x0CoasQcmiAJtBQAKDlX+2bnnAFIipYLE3nnTBVUkLF6ehsCqKHq9JbTgxklIsQYyQyAoGkIqVZT+tHvt/fBAGKWb19v/tNXf/wPzy8v/+b548fPtqub29tVCLy8uPDe361W/X5ngLN5t7hYGtp+sy0lr9d3oZTQdpdXl9st7zbbGIf13aqZL9g3V9eXTLjf7bbr6Bw753zT+abNaRj67Xq9QqLgG+8Dez9fzELhISYkN+uatpnNu9ZM97vdZnNjiC4sFpdXy+snppiHvn/zar26KTn5+ezy0aOLi4vgfd/vbl9+n1Np55e+9cjeN21MMQ6bfrfe77ZdN++Wl75t+/3u7vZmf7dp2+7y6mp+sciSdtuVZwy+e7XO/9ff//rXf3x1t4+fhuYHIKKmaZYXC+ZBJSNR1zU7x00TCCnGmHMmRBUB5sXF1c333+acTaY6WID1Q6o6OkJjtd133LYNEYW2822rq9s4xGXXVCce7xz8vKWzNb5U8z1yzkzoHIkIM7Yh1PhaymogplkkB2YCRKvWQ4BE1ZAoBNeGgAS1gmN98jtHZigiMQ2hCd2sY3ZStO9T9WUqRQGAmNghmEkpgEDM7PxsedUur3V+zV/f3m32uRyEkA+0wjgVVv6c78AZZ/x7wqn8uX7nlyLb7fbVy1e3q9WQEzIjEyBojdEiEBEYTg5jB2+v97auVfh82LOG4g/HVl85kXFKQIwqKjnLO1UCxjnMIckLUACyalQisAxKCozgpTABI3oGT+iJmkZDMAIjNCZgQs8cXKjFUQHFVMyUak0VAsKau0bcNDTf3saSyP3v/xv87d9+6qE/44wzzjjjHZwJ6DPOOOOMzwtD8OAGiKqmIjFGBPJNaJsZMQOClAKqqOrYEVYCmtQcYlOFtwgUApgBMQGYahmFJLXKk6GoiYqANrOuayA4dogMoAZqpiATL2eTKwJIkZRSSjHnosDV2VlKQe/NIMaBHTO7WmMw5TIuXCaX51KKc46d0yJjzT1ABBCReqK6YFG1Wm5GVUwBqiQZR1ffh7IMJ7IaMCBAYDZAdIxMIxNTMzCr4mYiZz27Wt59cng2mFZHtfJ73eCYK/FxqD825p+qjY7Yk4Z6Ip3HhHKccFT8VlIWqhgRpso/k7PsUXR8GM7JssNGxnm80BPRcW34KJgez3NQRx/USFOxocqG4xhrsAOTfSSgT/4c092PMmk1BR1tx6vIuRLQpqBaRe2l0nmTbBommh4m5vkQ+Pjg/WXHzjtmBjRAdM6BlBTzMGQVGS19tQACmAIYEXp2UoqqgavhgYTkrBQEpOCJSMzIOec9mFW/lNoFYtfNZt4HpE/GaqnaPpZ/+t13/+nZ8vll99//8rlK2m3X0dFiubh++lQQ9rthu1uLpKvLy8uLC+/CdrvdD0Of41wu5ouLy6sr5/xuu90PfRKZLy8uLy+ZqcS+72MsSZzDFtq2Y0KbrLcBTDSjqvPONzN2Xg08EaPEYStFhjgUwdDOQjdvm4ZBh6Ef9pvtalWQLp8+m10sL68vCUBSyjnt+2Tg5s0izJaINOy3282qH/b9MDhulsvrpplLLsN6nfseiReXV7NZV4btrt+ByWyx2Ef4/Xff/90//PrlzTrlT+aliYjMxM4xE9no2BKC49E2RxARiVQVAELTBO+996mkIsXMdrtdteepIY3pM6YqWhPG2TskGmJMKc1mM3LOu01owiexavkT8aEMgvrQJABCZHLBMauUIozgiINzqmo6UfDsCIHw8GQBYnaOnOdABGApD4hAhD44R4hoMQ4A4L1r2sDsEExyUgPn2YEDAFVx3vvg62OPnLt+/IxdSEWHrG82w/ff/+GbF2+yTCXLYCza+gBh8yjNPj7lTtJ2/vzO3O/HsVf3ZKEnrrtn/Ok48bZ6jy3VGR/G6ViNtZGZeNZ1pRQ/FezlsZwywJiGhXAIJd//8D3k2Vg/7oTVA+5kYmAGgFPBCHvvI+F+TpyBafXfyExiymCKIKCM4AiVUBiESCSnxETABI7IOSrEhYsjqr7PNY2jWlszk2OoJatd01BoYCh10vKrX/2UIT7jjDPOOONH4UxAn3HGGWd8XhCyMqKxazqypea9Ix98aELLzhMTmJkUK1Kr4U351FoTpwGQmRHIYMyEBlNAAzQ1FQM1NMDKF/rZ9XLLbdMeSFUDUzCESq2OQl0VURUVKaWoFEOQUnKRUgSJASDmwmrOweSzYDZ6Q49GgTmXoubEVAVqWT9iQqweggBABDJqsGnib6WuykWPmtiH4JCSCeMFTWpiM7A6EoaKhlop3QP7a4fzHKTCWtlMAqCpMiPagdw+sZyoXokHObPqWMHuKHY2MLQDAa3jugrs7YubeF0AOBLpo9b5dDl35JoB8WCaetrSKFY+2f/+1R39N04JaLN7K8hxGxwF8UdG2o471zXiweBZ1aTKSKXS0BMBfTTxODkJHtjnI8v91j1FZCJ2ZPU9MQ1jSpGcc4jsne6t5IIhOBMALCWrGiDVYnExJiARM2BC57q2Tf0emMl7BQOwtm2xit9zDk1L/KN8AD4CAxCDr1/e/ufffP2XT5fPH89/8fiy5N1+t0GHy8dP5o8eCd4O2/2w36+kPH32bH5xpRyy3pS4W928IuaL6yehnRWDOPQ559jvpAtFtQnsqMs5x5j3u41qds43zWy+WPZ93/e7mPapCHFpuiURaJZ+t91v1rlkIu/b+fzqC/QheCcxrvfb3eZORArQ/Mmzq+urrnUlDbv1SnICQO4uQlgsHj2bLZZxu37z4rvtZh2zkG8fXT1/+vgLiyXutxAHB3b17PnFo8eoaf3yxd1m1V0/MT978fLNf/7qD1/98fvdkD4hOWSgRUpOGT1679VsGCIxi4io+Ca0bVNV7ZJS2my6biYXF+sSpUgpZXW3cowcvEoRkWo4IaX0/T6mbACmmmMchoGZLy4uFMA5x8Sf7gr+VBjCuyzNmNqAxMyOAE1VhJkQkJAATZEAxgQT5x0jEAATOCbvyTlyjEQIpgbKPDo/MdU8kuKcC8E3TQCzUoqZIVIIHpHVoJTCntk7IjIDUVPukuBqu3t9t3252vzxdvf1y9us9x85h76fXsiUO3L4vRr52+H5MwF+1hz02/g5BDD+P4iTzKIzB/0uTmcUh0/NW6jbau1Q72ohkaMwwU7asUkxfS9u/l6ccNP1vFOUf3px6sxpDz+gP7i3hQiZyTtyhITGYIxGAITVQc5GMyHU+hwZCWYyQiA0BEVABmOsBUeQCBmBEHhyIiJCRDIzU/xf/+f/5v/4P//pxwz5GWecccYZPwVnAvqMM8444/MCGUHAN/P51ePGlmW5rOxwSdkFH0Jo28ZEtBQCGIvnVU6zSCXdmtBUVlpViMw5BLJa/k0UFMiFhtBA1dz89c4t50vnvAFMnhSjYTCOawEtJQEoMyJY1ZRIKSmVXESBiFmAVFGLVjpW1USFiNh5q4JYpCIqkgyUiBjZpBwNPkytVCEeOOcBUFREipkxESCLjuVuRh75IZhkvKoFkIDIBIFEiCpVPEqMEQFqSjiXXCrbXtcZiFgl44xMREBQnRkmysmgkiaVyEGk0boUcSTWlabajAed74FrODDvxzzycR13UAWPRPdRyjwRxu+uFQnJ7rE2Ryr8dHF5WOJN/Zz+vmd+MfLih11PTndyXjsehwcn65Heq4x0rSimh9Tat+j9WqLwcN0H/vk+hT5uySkNQ59zIgZPPvWbFKNz7i//8r8IRNvNZrPZ5JzNaplDkZJTyk9mc8dOU8kxEaFUV1pRjNF7H2PMsYcSEX3T+MVybkUCk8V+c7ca+r7K8z8VDGAz2O9f7/7+X795esGP/sf/6vGTJ87xPvYvX37HvlkuLj2F3d16t9vLd9/PLq+7xUX35Zc3r1/e3Lx6c/Mmii0Wl1dXV7uNy2kwlTev34BJ27RdN/POiUiSklKWos67ppkvF4tShmEoWlKMToyJXEql3w+qUHL2TXfZXSyvH7Pz2/Vqt7nLcZ/TsFhedPPF4urxbDbbr16v714N/U6KELnZ8urZsy9E9ObVd/1uvdmsNuttO1s+ffrsi+df9v0+Drv13Wq/u5vNF9fPHqnI+u7NZn0DYN43X7+5+39+9du/+8ffv75L6RPaPwNArVPJZAjOOULut3szUxUCC94V73IcpO0QlNCK6RBjKcLEJedHV1cx9m3bdm37pr0BgJxzTimnnHJpmgbNckpmxsze+T7nIeUY45+f3jrwMDgFnU4CPDUIiYTsGKv1uoqCqYqaIgAjApCaAFhw3hGSqWP0nkJwTFSt0QnBMc3nLaLFNNQHHhI3jW+agIgl5RwH773zznkyBANyTaNACth1s6I47NOrF3cvb9Zfv3j93evbl+vdTbGNaJk8509tgu5fGzBxLVo7CjOZnXM1wKAH2xTV6vIE958kPwA71no9bpmGEz+05XT7gRl/i8g7pT6nAz/S4IfOe9j41pvtB3r4A1veu/2jg3DY/sDh+gmj+sPD8t7WHrIznhg+vNXCT7i69x7+538I/BiM8RuiOmkRkTETa3p9ooIVK+9Ko52aqqopiCIRICFyncFVgviQjXB4rx7nOQeYIRgRjcpmVWYmxzZOFyblM1F9nFW1Nagpvv1tMc0mRrs4ZmqDW7RNC9CYOiBGQwSm8V9PGAgdo3ccvHOOmSvFjIzkiR0iIzBjnQsTG6KBCWnNtiATLiULgJH91dOLz3iHzjjjjDPOmHAmoM8444wzPi8QybUG5GfLZQNZnVYLvCJKzpP3hoSMjASiqlaKTrN8EwUziLkUKTlH0WImAGJQABQBxRCAvPcIBqrk4/buLsUBVBjgKITDaV4PUBcY7FzbdcvlcmZALuz6FHNJRVwIgJRTqscREVhdpBgSBe9VtYiUUoiImUVLJWeD84ykU6kZVQWorPdI79a8eOe4JOv7RIwgDyIV7JR+hVHjawdNnKrRYbFU1zZqiKoIOi4pq0kxEdclmaGJKYgpqioJytE0AgDGqzZVYyasboYHzw04/HMiZTaw0Wvk0MXJB2SUFB8FfHg4zUhFH+7KccH41tr45KSHBsd7el/2NB13b41ddzmIm61y/njEpMc+9mr8ZbTkIEQUAFMzPMiard7ew9L2/tE4iaBturh7A1wDCaaigIRIznlhV3Le3t7OZvMQuJt15P1yMXc5lziAChKmoq0gKVqxPKTF1TWD5X6XU4o5LpfLrmkBQA02m82b168ZEJrFzAccTaA/pQgaAMTg+9vtb1/c/vH1xT//5qv/+q//ZnZxaRvsN3dIvLx43HVzNF6vbmLMeruyLPPl8vHTL9rFMsU0DPHNyxeLxcViNitNs99vd7utlARIQBxCs7y8GlJMKZWSRKKW2LbtYjZvgo8pIoIW6/NQDF278L4BpKZpF8ulZy1p2/fbmLNrZtePHofQtE3rQPubl3cvvy05kXOzy6vFxbV3LjiIZS/xZrtZReOLZ18+fvrF1eVlSX3c3sS+B4DF1ZPrR1dlv9ps77a7vTXd9fWTocDX377+x19//S9/eJXk03M2huhCMEgxZc/Wtu3ru9vZfAZgZRhy35e4yzGAlDY0kgsgoOPQNvPFXLXEvk9DRCL2QURyzgDQNG3SPTuXSzbg+ax7rfbt998ZOREldvaji6N+TrxPBD3CQFXRRusKMLDqg29mJszonONK0JBzDh2jQwATBOvalgjATLQgWvVkd4yA4J0jQlX13rdNg1SdjlgBjRy50Me87dOL1au7ze7NavdmPay2w92u36e0L1oU9BD7HLv5QdhBfokgINVN5fDEPHDQdvIU/cAoHeNzP7Dnu9s/IBS19756+ufDTwHvo0F/oIV3T/SjJNUf2v9Djby7/SFb/pQDP4r3jsx7qeGHDM579/nhLT8uNP6zgZkpKBzJdDhUNZ52GYt3VOYZAbx3aorMVoPj4xf39JkcI8p4yBF7Tx0FFUQgZjtY7Y/ZaYZYywAf4u1TyP103vPWJUxTCARAsOqh5AA8UkB0BMRAjJWADhMB7Rw5rhw0OSYm8kSBmY8EdJ30EhESYfDsnOPgqJtrs7j74zcmqA+NcJ1xxhlnnPEn4UxAn3HGGWd8ZiCqOGYAMEQF05JTjqmkDABmUogYkQyllJJLNcMAMOdcVbflXHJKuSSDSv8m1QIwilYAyDlHpqDKIe3Wey2ZVPkwxZ+WDxNTaIbGTCGE5WKhgOSb0JSUS1ZFZjPIKYuKmXnmygOM+hpircUKc3Hee+9yKSWnUnLXtMxcU7YBAECr0karRzShaAFTZjf0WdXYEWZ8qPq5ctB1MVVzzWsVRQRAqprlWsZ9lNsgAEDVPRNRFQMdfKK5Vng3nfjj48LooCy2qtFRRASZSsNX0h9gqux+6BJMMuPxeDshjSv9e4+OPVwVHM6NOFqHnFDhR+Ydj9x3Zd8nqfJ07HQR+NY5KgE9Lh5tdAmpZDpUR26kUw4cAAwnzRLg6N5KRjqakpz2fDrbkSIbR2lin0+v8N7QAowWHI4diWgVXReRGFPOGcFMpe93pSTLlIdeSmm7TgHN+bGAkEE/DBei6BgLKSgRmqoUsdCIKABWaRZ0rYHxaKf+KVeZBrDd529e7f7127v/8GR++fLm+ZNHFxdLsrzd7rZ369nispvPCHHY79Iw7DcbVZ1dXXXdLPgGDbdp02+3ZOqC9963bSvFkXNimkoOjM6xCEm2IkmllJLn83nbdCG0+35QLSLqfLi8ftzN5uyCquScVm9eIlEpKbTNxeXVYrGIfZ9i36ch7Tf7zR2zny+vlldP2vk87dbru02J2xy3qmVx9eTRsy9nbWMl5WFb0oBgs/m8mc1DG+5uv91s18Z+trjuLq6//s0fv/r997/+w8vXq71+cr7GwFRTzkmLlmhOG+8qj2yi5CwP0TN7x6CahpjS0QAEkWKKqlKKElM367z3zjEgqkr9SPgQksAw9EWKGagBEDsfPvFVfDYYgJpxLRLL5Gq4bHQoguC4bRyzeQbv0FfnDTAzZca28YioWkQLIjZNcITEUM3xEQHNvPdNaNVQAASxGIqRFljt8+ub9fevbl/drN7cbtY76bMWM3RszI6RioDKW119T//N0CZuCsDMRNVUx2yVKa3Epp0fMCKf7B34MxTA4n3ribeUvD/DDn9a2Emlu/e++tFjH36iH925nw3qN/xoFwan84mRiaZqpV+/+plCCICITDrF2Ef2eYz5jGzwD42eMYJVX/5DuAhPC2MAAKBNkxtCMEBV/QFXj/GYsedAiAzomDwRM5CDWjQxIHpGx8BEjtE5Dt55x47IM3lmh8BYXeUMwJxjduSYmuB88By8my9Ls2hehH0s9O/4tp9xxhln/HvCmYA+44wzzvi8MIWCWoa0ef2qz+u4ed3voxYl5lLEwNrgHTEDSimllFyySGGG2awFs5jS6vZWRJi5aTwSlJJqYT8gInbMTivvoODFo8qsaRrPPNYmB4sAACAASURBVNob13/HEuQGYAgGoCpo0gSfipSSHTOiIymqZqDkMGctIs4hICoAjwJSUzREAwDvIXgEMzQkYu+ZEE1ATMe5PjMz5aIIwOzU0NQMIATXNt47SoTydiH0Dw8jjusnICRiYB4NN4gQ60hQtbOo1cmc41rUEQCYHSIVEQQbyw/WEcDRs+NEjjMJlyubYQdnZ5jysU945lNZ9uSucSIGxrECIsCoqZr2g3EhPW4c82drX8wqOV5No6kuGfFUhDS1Mqal35OHv01Awwm/A1B9NE5HFAB0vEY9/DgknlstI6aiIioyZuxWQaIdmHMwG8u7wUE6WoXSE3d0tB0xG+l5HGvK1aGp7gFg5hxXSxIRGfp9jEPbtciO2DkgMAE0ZHKOvQ99ygrgfKiDVUpOKcpoZYPExPUWmPkQqhbroe+2ByMLvFoN//L13f/w138xf3k7D/zF46vLy6ucdbPbGYC7uOraNrDbAu37YbPdCehisfC+mc86MBuGYbfbhBxCCIvZjJ0Xk5RjykPKfdu0ngmakDNIkZgz7PcGEHxAJO/bIuhDmDXBMRJqn4ftZjMMfTtf+NAuLy+XyyWC5n67226kJFSh0Pima7o5O06p39y92azeqGQkmi+urp4+W1xeatwP27vc7w3Qt23bzX0IMe5Xd3eisphfzubLfZ9++/Wrf/zNt7//7qZP8unlz2CiOsSYfQYpBBiIHY+VpTwHMgyuaZuOncs5qSrVMJFoTmm/2xcRTwwAnh07x64WNKT6lHA+CFqMUUS6blaACMk+yot8VvzYk5sxU3BN61zjufEEImjKhG3jutY7NkJFlMazc+hosiMiJSRmx4Yh+PmiyzGK5EoiEWEIgZiLWVZLAkPRKLAb8uvV7vs3ty9v7nZD3g15GDIYARGIMjH54DynIW1L/05f384/UFMwYObqxYFjJbSRqVI1gHLQRD9oYN7nzPCn4NO29vCm8PBdcLLllEV9t51Degce6gccA9B/Kk4/2qetvW1bAQfe86ON/RTS/Ad45J+g7/6QJv3kcv6t8VYs4S3R98mf9dV7B+IUiD4J2Yxh4Gn/EY7dfDFLKbZNyLll54BQDXSaWBzj6YYf/fAhKNa6zWaH2ddxbKcJDwKNEwxQKYUQS47vWGLZ/dMhAiHQNCtjREIgMDU1AzQCMzRDMAQjUzIlMzJDEQApSkAIXEXhYArKhkWxaHYlUfJURDpJkg8zlDPOOOOMMz43zgT0GWecccZnhmkwK1agJNbSEJBnc8zscylq6pm5Vo8iNoeibCBEEIIDsOCR4EJEkLAmRyMYjDo3QOIq8AA1UAuzq2jy6Hro2oYI7nlcnOhUAayUMgxxv9/3McWiyN4MihQiNrOcc9Uyq2QAUDXnHBFVs9G6jpBSUow558oRaFEEFBEzNTBMwMxEJDKtT1RqZmtOGmNUlWoQ8iNQ1yNIRoiINcOzyngnK4q6/CYiqvXEqu6ViA/sMCEQMwBURWzV0k5a5bGpapWISKOcZ1qTTQOJNhks1mXa0cTiRIEJOHEBI4F91BHZJHA+0TKf5KSOCia7t6w8sOKH8oJjNGEsvDid/FRBjTCd4CCgpsMpzSa+fGSc9ZR+PpDtY5lJq2MyNj2d6YT5Pr1PdtTaf+hOAphZKZJznjOJqUghpq5tmiZIEXYuNA0iYmhml95S+fb77+ZNtGFP3nFwLoTGkMkBEjpW0ZxzyUVyoVJUJQ77tmnYDDabbj4DRBH9HJzCep9+883qq292j8L85vVNQHny7BfLK8zlVR52dznNmuV8cdldXKvbD7tN3NyyRFxc+aa7uLyYLbq7mzex31nJF5dXFxcXMSfdSd9v07AHyYvFRZjPs8x2ux2qxBzz3aoJjQtN0y4AWaX0d7fD0GfJxczI+XZOHC6urufzGUjerl7vVjf9kHzTdMsr9i6ExtS2qxtJw27zZrNaCfDl9dMvnv9Vt5jnfiP9TmO/3+3axVVo585xSfv17ev9UObLi9nskox+/4dvf/Xrb//pd9+/vNl88lGdSJT6YySeYkxtM1vOL9tuweSbZgbGRMGH1rWtMe/viJEIoKQsuRQR33hmznGrIirqfVgsluvdXopIKYS+bTpT9cEzOiRKKX3ya/kEwMND4/izhtMY2RNWn9OcM5t6wsb7JnDwFDwRKhg6BkdAZMxU/dOBkByTAYCllMwUkZBQTEWr07+pSRbcR1nvhtW2v1nvX9xuV9vddojFKBcryo4YmRiVXSDnARExHzpuUwDq/Vc1xfVqusmowazPnsnR6H5Y72Pj9ElZpE/b2kPav/9QxffvfMza+YFmP/Bs/kl4K5nlPV063fagxo57HdjVj/LRH7wdh4H5Mdf6Xm56irxOXZq6+PBm/3Tc69jBBON0bnH/9cM0AYlMDVGn4MWoXwZQmHwvavHSpmnYcRHJJedcgNAAbZyE2DSvgTEvBICm4LeavTMaRmCVgFYdpwtjetgUWTcDHQ2aDBFUREqxD34b22ECYwI5lQiGBkLkCB0ie3AOmVDJhNAzCZM6spohWJBpJKoZjQmmxCd1juvXgyMiR+QcpqTZpAhSsIc+Y84444wzzviTcCagzzjjjDM+LxhAAJnRIbbeEbbQVms7FtMxWbIWchlJSzQ0Q4VREGZX19cy1WIiQl/FyFg558pGo5mCqm8fRZDrq9i0zdF2w6D6MB8cHgykSBnisF6vt33fZwFyAGiqITQA2Pc9IBAhRDA1VfPeA4JIMTgaHJtBKRkMiPjgOVFPKaJIyIQqI09qqgZGRKVYHNKJWccpPrzCxON66j4LU2XApmpA43Ksss710PqLVRuNamRca59XumUaExwrqlcfD0QEZKbRXrqWd6+6XYRqqHyga+EwHm+tC+sQjdWARib5tCrh25d4lDtR/fsoy5kOBDOAGgM4rENxen00+hhdVceTTi0jwehVMl7t/WNPoCP9M/JCKqRQZc4i9SZMb6T7Orv7GvCDjPp9MFFLOeeciHjWdim1cbPp93sKQVVKySklU/A+UBYwFbP9bj9bPgI1YFbnt7udsa/e3qagpajIKCk3Q9CmaRw7I4bFfPXb3+aYPgedZABZ4XaX/+5fvv6bZ//lBW8t7sHC0y+etV/67Xq9Xm/v7jaGfnZ51XRdmje72xfb7WZI0i0vFxcX19eXKQ45591+G1Pcxb7tOgLtGu+xjbFflezbRdMtl5fXpaR+t0nD0A8pGBANTGRim+06xr4Uabru8uri+tnz0M5KzqvXL4bdjkHMoJt1y8ur5dX1kEtMQ469pqHEfr3eZLGrx0+ePv+Ldra4efXCJGtJkjP5ENrONyHH/erNq9c3r6+++HJ+cRVj+ubrF9+v5J9//+LbN7s+P5zZP2VS4OTz/p4GDAAR2qYNlLlkR8RTcc6Sc9RStXub7eZiv3/25BkCxn4Y+qEJoeladAwZTMSInPeVDEk5b3cbxzjvOokxa3bOlSIOsV0ul8ulqvxMmYj7HDSgIQETeQRPiKCiJefYMASu9kjGbOyQkcCI0aB+XQACsIFCrToIpCLb7daH4J1Hdiolqw7JREsWigXW2+HN7frlzerV7eZmE4uZEQGRAREToB+TUrxH5qJHL3A73tf3fPTqE8PMRGWMRU6hRJgeQQe2C98pAPhx/ew9se4HdrkvMn1r+9unOHnzngYcD4Vkf8ITBk9U2wde9uOtfOxEB/L0o009hPl9SDv1qwfGr7kfbnAcW5xk3R/loN8a2PeM8wc46BM580PU2XDoGBxo8h+r0/6ROL2Wk94CnHyzTn+dvPnGTuE0J4HJl0zfabBOFg6hbiAmxw4MUor9MMSUkRCJYay6bNM3eA1BARwJaBPRtx+PZgjGRHogoG2U8E/FnNEMUsyASITMZKaaR8P39+H4+NCiSROqiqpDYARGDI3zDpnAM3gCT+S9K56LCFPVJBghcJU/ExADgqGNsTckcIzETN5hFlRX1MzhoUbKGWecccYZnxVnAvqMM8444/MCgVoAsUqIckrCWCuBCwAgmOhYOYqIAA0UsoiYGI117bxriNiQck5gwijsmIgRWRRFAYlMUcU2cX97J7lgKpgKHNYKpiOhaQBqmnMBACQaYtz1w5AliakhIXkvRCxF2TEblVKKiKq4bIhQjaGr1AUO6yUEBKkrz3oBZqaqxMTMUkRVTJWJKo9pCkXUAAGqSBvvjdaHRtEA1MzEVJEZjJABTUHJxmEDk9GoQ8xMtf7OhSvDKkUck3OupISISAyW6ylrGICJ64INR+4fiAkBVUc/64mqPngsTrQyjIMx/jkK1CbpMSFMIuuJdJl00RPlcF8BPabOnvyHh6Xw2PrIrk9rRTjWTbMpf3bs67FPI1cPxwWsHQ5RM1U96pTMxkRXNTOFkZUeifUPLfKn7r+90Q7ngZHARgSqdpRIKe5LzkzYhBDHRSmBoYiWJNpZ3u/265UjJN9gd5Ek7+7WzpEiShyG9aaUvFguh+3Wz2ZhNteUYj+UnEE0pxQMpJSDacgnhwHsc/nq65dfffvk+eLxY6Q3X3+j/XD59Gm7vCoY7tJqdbeOIovl3HsfFlfJXCopb1a5JITHnt1ssRi8zzlvN6s4bL1zznFoWvatGhIzaEbj4ANfXKUQh74XES0ZEdUEnHfEV7P5YrHoZjPHGPd3+32/2+5zKW3XLi4ftU1DTP1us9tvh9h7R4RQTAv4R0+/vHr8tG1nOcbtzRvHSCFwt5h3HYJt1ze7zSYOaXnx+MmTL/uc13e3L1+tfv398M+/e/FmvXsA/XxgT95Wz33sMETE+h5EJmZOKQ5x35bOkIe4LdK35Mxy7PdI7KqbEaESuuA5UhlSGWJMOcYICEOMpRRELCURISMVKcyUcqI4mArzwTz/KDn8ke+IzwiZvjaQkBwGZA/AoGBqWgiLc+SDsRcgFNOYEiMwATIRmprWQJQCmKpJ8c4DkQGrcTZGIcE2M+yHstnGu/Vwt+5X693qbj3knIsy8RgXGy31GdADsiEBkhgWAIG3/FRtClvd3zoZAr0r+YTTJ8Y7HOBDKcEH7PWhpt6/3U53ON38/n4+BIdDRprwwYd95PUf34EHN/iBsLF9ZBDwfa+e/vkDPRkji3DyRfhu/8Y3zj1PqrdP94CBeWCXPhXsxFfknd7C+OS8/3GAaYIwBfvH3xXHEtDvBCjqXypa6yfAEPuYepGSU0oxIzPyu28/g9HHA/RoGmZvaaArxV1kNNbX45eBoYBMFLiCIqAZqaqpmh2y807bOm4gABARs2yApgamhITACBJLykBgniEwNs7FnJgoeHaOmIgJHFNwDtGIgBWYkLHG4JkIDU2RFChwYB9gUHt7FnPGGWecccbnwpmAPuOMM8743GAFQ9F93wuUuN63IRCRlFqEsFKyBmA0FseDXLKYAhMgErF3SMQIULKYCoFxViIB5FJAtXpKqIpEsf2+pBi1yDiPHz0l7HTNoqpgVv2FvQ/oALKIGgKz84iEWP0zyICAxNSYq9HHSEAzjKulWs4G6i+1bNS0bqkm0MJSlxx4XM8giQ798FCK57gymLwdBA0EamZ+JfYrtVu52YkkrWpftLE0mZmpsopo5dqJqygbEasYx7Gryz0iMgAVZWYkVFUmJiar9OgkPzpkmMJENI9U70QaTxKqaRMiTN2c6OfD9b9fCmrTGvRA++LkM1JfnkRS90ds4rZPfUNHo+aReLbDqepy0szUxjs1maxUP1hTFRWtUij8mPzwgSv2qtuqqPEKQnSOi6CIIqL3wTlvgICkppITmDE5dB7FPHPTBDEaLVacNzHPngBBFZGapk2+0VxKyijahNY5j/i2C+2nQhF7vR3+/rff//Lp8svLR8H6m5evXDdbPH4yX17mpLvNbr/bmpbFxbKZXSi63e4uDrvt9g4BvQ/Oh845l1MZ9iVHKalpmjYsfNeNrpk5l5zItaFt23bmnZeStcScC3u/vLgg4ovlBQLklPb7bSqx3/ci6pt2Nps570sRiUMpg5YBSwTgrFBEL66fPnr6C+9dHPq431nJhuycb+cLF/x29Wa/25RS2vny6ukXotDv+k2fXq2H//irf/369V0fy+ciaQxEVUTZVzOd+lRCMyVGDu72pjcURDUTKcU3jIDOMzunYEAopYAIIVQLo1JLGqasWnKKRIhGOeX6cMs555Tos71JHnjJH6W7EYEm6yHH5EBJgQiRyIia1oXWMRuS1FQNBSRDMUNA5xwSGRgSARFULydkdmTks1JKtstpM6TVene3Htbr2Pd5H2M/ZKj+654IRjWpIRuwAopBURMpBSxCiVJOzZ8+dEWn3OuR/vm3tTv4eeFepO7TNfWTmbUH9gNP9run0v8RjX38i8NgTPT54Pvp8P9P8xb6N2CfDyf6MP1pcPDKemv7yMUfXjK7tyce9pqSCgwAnGPvXc4pxlhKVjNAZGI7aKTfPgvAFHeuUXnEez2pkxqTKThPiABIbz9FiWoQfwwjTBMXe+e6EAAIjAGY0DM1RA2AR3BMTMAIjpEQyMwzBqbGMRESQeOdc9VRHrzj4B2CEZlzxIRMWAuTOEfEgExAHOZLaBduEP3zPvbPOOOMM/7/hDMBfcYZZ5zxebGFRQsRdf9mtWaNZX23XMwIIfY7ETEAQjQARauzc1NIpRiA896H1nmfYhnpTTMYq64UMxAzFTBF4sqCWoGQcx76HZTsAQjGonullLd6ZWaI0HWN7zpyTZ9zLqoCiAyAqvKWiKauKGoZOkR0zqmqiNBoZ0HOsZkNMSKO+lwmrrXRawspRZVSWcec83a7rj6jDx3Heyy0gpRJk1tfRSACJJgkyYhIzAYqOdU/HbssmsxUBBHZuco7jwS0mfO+GpCyc2AgIkxciR4hoTKWbj9kjtd148gHVe4Z71WCUhvNotGmVNkDCT1eyrSCnHBgmMfrrDW4xhMdSW6gWq7QJvL7IMQ+HTCESdx9MMQ4nOY4mFNfdHKBRjQcS4QdnTimLOlRRwnH9fkhUdgm9fT0FrvfnxNG5CCGrKELNMLxQwBmqlArSwIxe3SOnCPnDIARUYpD6Lqum81iEu9d6DoyWL987dhhztL3PJ83TbtDNhQEsxybEJj58ylZDSAJ/NMfXv/VF4/+8umjv332aPPqm83dLYXQLS4urq6apl3d3vZ9BKLLa+89dW0AyDnG3X7TdTMfGufYd4153u8xxjTkgrm0HrxzxUxlSDGCEwToulk7myHY6va1lOKcW3TBu8Bkm816vV4XVXKEak1wXdc0joZh1/eRENuGZ8H3mlNOKRtQePr8+aybDdvNdvVm6HfM7Nuu6zrvKPb73Watot3iYnH1ZHZ59fVvf73b9+t9/sNN/x9/9bu7XfyY/PnAibwrr/sI1LSUoqrMzMBqlnPmEc6xK1LGVAMkdJxzUVVCcswIICoxRQfAIQCi856cJ3aGaFJyiuPHGbANDQLknEsRpkM/8QGd/Ohb6sdzWD/IQRMAI1aZ9phUboZmwbNDMLNu1rSB0QqiIRox1MQNEWFybdvWWqLEhMSELIpIzoUgQCnpatd/9/r2u9e3L29Wu10uCXxo2XvfLupzQ0nNDA1qRFEBslgUGZIkLUlLgpJgNPj/5DrcER8kys74pPjJo/qZbscUMf08rf858YH3/3up5+NB93cDeI+LRJ1umFm1Zsamadq2EckpxZwzEYXAITQ6yiDeat+m7/0x6lyqz9XpCUb9wegRVicp9BYBbWCiNWqmpoaGQFreubSJTEcAB9Awz9r2sg0tUSAMnl3lkZkcIiN4Is8UmKrRcxMmAhrBOfLeISiheUfMY8DbOXKevWdiBudcu8jcNP1Q8rve1mecccYZZ3wWnAnoM84444zPiwTNa3j6S79u/OyiewSXi1njCST2exUxq7a8ZmDAhACmVnIBwOBbFUkp9fu9SAZTQkMwOqhODGoNPckqUqSUYkEGngUIjGPtcDvRrsLRRpQAPPPlYpFEMqDzrSiqqBrq0QFYRZUQa9U+VVVGRDdKcomJgmM2s5ILEpha48kH570f91etRW+cc32PJefqwpcdz7q2pJjkbWb8/ewL3t+MBMhAQETIhLWiIHN1cKZJhjymo/pQqWGeyg6qKCISY6WwkUZpcxVC2iRvpnuJ4eNq7EQCPJldABBBXXnZuOADALSRkq05q6fy6CNZjFPLWBXKo7MzElWXDmCrQQcbD0OqFHtVMx/HZiKtq7nGCa89smijFzQcxdMnHcCp2iAqmpmhmYGijeMDk/x60i/VAmHv8Mv32Odj4ycv48EZRBVqgUfHDApjuSOTmCJ7V5Ls9v1u17uxPCeR8yE0jICxV1Az62aLmDc63hCcdV3abrS2m+IwDKvVbdc0wfnc9ymlUop+lhqE0/UBvNqk//urF88fX//yL/7b9vpis7lJebh68vz66ZdX178g19y+ed3vdlD2xBrabrmYx8bv93uzVHIxdSG0LoSFf0R9v9vvV+tdV3Qxm6EhIoemQQSToSRwPHO+8aEpUtC07DboeL3f3G22USEsrp1rry+XjXclx+3qZb9P5NrF9dXlxcJKv9ts+30GDsuLi+ViHvvdsH4V1zdZxObX3eWjNnDabzc3N2lIzWy5fPTF7PJ6dfN69eb7bO77m/3f//bl716uo/wwG4Tv/PLuS/BDfNVkEVuLTA77XkshZlXd73spIAJIzofW++b1m9cIAKKSCxGXImKCgEVFVMFg1s0uL68uLy53a8k5pzi4NswX87xcDjEqCiLUKNSnw/szGz6CKbKDh3KeUzMK1bwZmxBCCH2/L1ZagsCOPDE2Jcs+Z0LtuqYJ3jEQISM4ZmauBWIRiIkNUNQMOA5l1/e7vqz3abXpbze79X4o6sghmYKj+iQrZgJmigomZsW0GBSDbZahSLYxdmSExVDuW/x8YpyZoh+Fzz1cH2n/XpzyjAfjISOG975k4cjhTv8zPMm1MrNSciklhNC2bQiNGimgc+F9WgCrcXY4hMwN1N5j3FwnNKqTpc40LzppyWz6qjYTFVLEkhPIey65TnEJIDCHGmCTAqqi1ZoLgB0QQS0xQlQYjdAxCXhUQiZAACEURlRC+3/Ze5MlSZIkS4wXEV1sc/fYsrO6pqq60SBgABwGRDjgio9A/wI+A0P4EtznMt8AAhEOALp6X2rvrtwqY3G3RRdZmBkHUTM3XyIyMisip6ahLzMizExFVUXFVMVEnjx+DELGyETMZMYGbMBmDKbUgPeOkRhNce5WZsyYMeP7wExAz5gxY8bHxQ42f8z/UqNfrOqLy0uMTe0QNTdtq2pghliMNwyZyxhfkoBC5ao4hhEHFM2ZTBKiESiawtHHobCakk3AxECJgWvh6mJdtzX1SeV2MoD3FH0E4B1nFU0JXcVUTJa15OBTUwUxzcDMTJIL7aAlklJVEYqmhMxELRXyElAAqGRdNxORTESIJgKq2UynCNoSUMn02OT1/WaqhYwlLPJvImJmRLrNCQ+gxQaaikgZAZCJiNCocDDFeQNLAncwK/S0GagpIjlmLaqg4mECd+JkJ2qoGCJOcaV4m/jveCFGRxH0Ge08yaCng5TY1qN0+oxMPuq9pqSFZa9Cr59sqk/k8kn3Xao68d52FpZ7W/nbehxnfGZgZcHgTO5saqf0WkcLkEkCfeL4b7+Q+76QJyuScxwnw6f5rIgggeScYgKDtlkRe2L0vvLelylhSGkIoapr7xiZQPI49p9/8cVqvUFVScm8Tzl+/fXvnj59evH8KbV101RXV5cmIgjN+jJ9tk/5HVmPPgyywW9fb3/6iy/+7U8++Z/++/+yff1lt7t5/fLrQx+eP/901S7qFy922zc3298xY1Ko66b2tVXCiCI5xBCGEV3t2qZqF75ux3GIId7cbL3zlfcmgmgmOOYcxtH5um2buvI5xr7v9rtrIvB1s7l4cvH0E1fVse+212+67mAGdV2vNsu29jGMu+vrIcS6blaby9Xmcjwcut22OxyySNU0q6vLLHl7sx921/vt3vzq6eVTrtub7W67vW7q9s1N+Iff/O6v/ulfgsAHovQf1xojIjn23se0Dd0OFF1VRU1VVTvn0xjXm4uXX32ByKp26A5m1jRN6PbDMIDZerHMi1XtXeV9fP1qGMJiZc5555gYnWczIyTn/as3bwguLp48r6uq6w4fJ/T+ffTUd2HTM3SHT5qeISupQ1NKhArsDMysdGVqAAZEyN4xwGSF77wnJM0qOi3gZbEQJYruuvBm2+32YdfFfR/7mJMaeY9E6AQQy0+OIGTDrJpMs2k0SWZR4ZBSKD3p1Mnht9I+z/hXjflG+G54r1HQAzeSe73Fw00Gx3FbkSqzYzScbMvu9XvHUc1tdRDIHrGqKKJnAAFVJCzeXffLHNfzy4DEHnpvwDEThmmRchMRI6IqgBrqNBCaBh2MWPQYZiU1MgGYTJlWCUFLR6hKZkIGVNIIlKgNkxLeBVlEUjYCI5v55xkzZsz4fjAT0DNmzJjxcfHnf/7nP/2P/5syLptq0TZAmdAQnPMVFAsEkyJxLSypqWrKkBUVucbGV1dXl6aiOZkm0FwS8RVMdKUZITomrDcjtNcD//CH/3D1M3e4TjHfStHuWC+Yicg4jod+OIwRmAHJFEqIpWMWsywiIt451TrnnCWrKhGXdIKFrkRCBSsuyYX9HOJQpjlqpiJHP2UxVQRkZkQUkSTyLQb894qeLCfU1LIBKpGKUUm7flYAEVEA0EQMVIWIC3tOQEwqBpPw2exIQJezEZng5IDhnCtzN3aTRNpMywSuvLnHteJZLU8ydDjqkY/C4EIhn+TJJ+Icbw9156qPemekSUc9BcjaUdl8VCcfKaqT1wYeT1Aqh9PZjzkRp2T3qioTB60qMp1TDWhKLHSrxSTEQocXR85JaX4k6M8Y+OPF2JGpP95703EAiVmyMjvvmxSjGcYxgoH3rm1rUAXNjsl713eDgoFjf46ncgAAIABJREFUZMfeVZUvdDmaac5D36/X66Zpij+A8z7GYKJLRKq8d46PZuUfDwZwGNMvv3zzf/3tb374fPOTp1dXVdvtD8PhsIWv0mK5WC6fPLvyq2q738cx5C54l5zDyjtlUjU1Dln6fVfX0i7azXLdwSGGqDlHldq7tmmJKMQ4DKPkjKbOu6wSsoCrm2W7ubxcrtaOIYeu273pDh1w9ezFD+q2zcPhcPMmpgDsiP16c7nZXCLgq5cvx2EE4OXls/Xlhpzb7behO+SYsF780Y/+zLWL/aHb769BErebX//jr/72F1988Wr3Tvb53h38Xmq+u7sAGKjaGMKalInZMRP1Wbp+WGyuFuuLvh8MgJ1zjs2AmcGxcw4Ac4zOOSIOMWRJVVUz8/QMGAzD4L2vKg+oMYYYY900dVOz6088yWN1vt8NvcdFnZd+hIN+3z7wvJxaTnnoh76uKgRfVYu2Bo1ZMhq2TVV7h6h17YhoGAKAVq74djhVyAIGqOzGmHddenPTvdl2N7uuH2SMmgwVCMgBMBBhMXpSBUZgFrPDEKPkBBpUo1k0y2Z6jJw/Pupw68gz418b3mfN+A/2q/9WPdIfOh6QzY/QuohITCq5xGHVdVXXtYiEGEIMWQCADCCL6v0H1u5bcICJ6sPnGhEdcUlYTfzI7yzabQxb1iw5a8oPSWpCImKTdPQLAzNQMEWbLoPQMZaIuso5z+AQyMw58o6dd8zkGEtcHHNxRwPHWAyHiu8QIGmJqQHIYQwhS9bvskA4Y8aMGTO+E2YCesaMGTM+PrKBaR76DikeXnsi77iqalGRLKppcpBgIiYmNgVTIwByjOiIyAgAwXIqXKaJWBZNuUwQ0AxMEUwEU87jkMMYQ5SkUNS353UxAFHLaiFrN6b9EA9jtOKeDFToRREVlayFQ84pW3F/VlV2ysSAKCIiGZAmshNSEa1MzPjRCGIyICxuywCFIzazMcY8jfvv4ZFI0PuzA1UAsULvTmJwVTW7S4DyZMpRvB8MwEjNyKx4v4qYGiLYRIXfCpyLBjkXZTRATqnMuSilW2cPACS8MwV8MO165JqONPJx44O53HR6OAmfb499R0A9FTgeDM9Pd9RKnimdb09wEiffapvslrFWALPpexdVVZnSTt5BUXSbAWKRVt9mUTp9BXg671T3IzM+Ne+UkwhJ1QCJiNUwJQWjsnJAYIgGJgSKACGFfbf36aJ2VJSew9CLCKpaFmKu69p7V4hxA8uSUQHMUKVyznvHDzIjfXBkga9vup/+7LM//fRJ89/+mx8+aS8u2CPm2HdpNEtLd1W3yw1Vsohjdxi7HSolUyLyzrNvKEvfjykENGibZr1cSSMpxZwTIgJxVdXsPCJKlpRCloRE1WJx8eyZr3xdVWZ22G5D6MMYvONmtVldPBGRrjv022skWF48vVhfLtuVGex3u+HQmcFivVpuNr6uhm4X+l2MkV19sXnSri/6MfSHfRgOdVV/dTP+7a+++vlvX3ZDemdLnN/YvwfXoxZDhBarunLkELDcMCXXaYhJxXJKotJWHhH2N9kQvHdlMcVMh2FEhMVi7b1HBBHJOQFAsbAIouM4MFNVVWaaUnpLJq7TnXxOYH0Lb4G3FfoWtEe5eJtI3vIOAVU1xOBRHQMRgYGpMZOKhZizGiEpOqAKyCNSTKkbY3e9PYzx0IXdfuiHOEbLmXIxDppWwQwQjFlUk4GIZtGgucsxqmawbCZmd5INHqmpmcj5V433oZu/W5mPjrOfwkfO/oe0ZPI+zfVo53FebGJxj6mhAcCcc+z40HX7/WEYggICMJLIHQLapqVpsCnr43HIoaanyKlTmBUiCmYtKS9Oa/MTe12GXtP4Eo7ObPqYH5Ydl7oVIAGMkvsAarlC8whM6IgcITM5opq5YvQEROgIS0QdETAhERIWlw4gNGZzTEwlpzcyI5Ehk7LjlQjXEQjZzXkIZ8yYMeP7wUxAz5gxY8ZHh8XE6g6yT13f37x0hHVVLRarlGJKUUTYMTlXIiKZnWZBMEfsvXfOqagyAROIIAASg5BllVFzFpWSuk0052TjIeGbEfe7PgTJAmJ4x3ujZI5Sy2JJNWYdkw5JFay4IjMSIxqImomZqgEIxFsWkhWZAQBFJIsimQEUt2gAKFkHVcVUJ/0JTKnsjtM7YSIDS0lEHyWgH/NJuJdcx3QS/h4TD5Yi53sioKkeswJOlDEhGtLEIB9DLo+T0jsTouMk6wHOAlLPNMVnO5/2Oqp4jkUAAG2yUMSH88RJzYzH98fPSoEzeve459HZ4x7VeybEfmAQCcejw70Np30MYIruL1roI+E8VeXEP0/CKACYnKvP4nePVboVZd+2yfQvTSkZwUyJSJEEUBRUjNkhgInGEIkBEVQl5ZRy7sdhE0KNlar1fa+AItlU0Wy5XI77nagCohHFEIo7CxlACCVE4GMKoMstgAbQjelXX735v//xs2crv3LPPr1s26cXh/22H8au2ybNvlkt1xf1xaZr61cScxxyio4Ja2P2i6ZF4K4f+r5PIbx48bz2Xus65hRC6IcRgRaLtm3acRyHcYgpeub1ZnP59GkM49gP3eHQ7XeE0C7atl1U7ULjuNvt9rsdmq7aVVvXi6urFPJ2e7PfHXxVV3W9WC3Y4WF/c9i+iXFkVy83m/XlVd/t+36QFBixj/rTf/rtX//i8y9f798if37Iibx/oz8qOgbJgogl62CJQqgqD6ZD18WYzGwYhxjCZd2YwTAMOeemaVQkhXBaBWPviVnVYogxxsr7EkSSkoZx9N4B2DiOwzC8n0/Lvaf3G67x3Zvfm4MuSU6NDAEMCZmJlFQlhORqR8TMZKoqgORUwRCIHBEDeUWnxinatkuvt/2rbbcfUx9yHLOoITKU9UczJAMCI1NAMYpgwTSKBsmj5kEkg+mDHIOnPvQPh8Ob8YeNb35wPgLedUb8g5bt32uud1zInfGMmZUMhKWjYXbO+RDTMIZxDIYESMXF6NilG4AhlR/3B4JxK+ksjuM6ve/iDDDZdB1HC2pnOTAQoQTwFbv4ew2uZgjTkpYAxCyDapZcgXmEomt2SEzgiDxhzVQxOUYmcjwJKEpCQkIgRGYgAkTxzI5JVBHBlR6R2VxVcVJnWrfKjh44Us+YMWPGjI+BmYCeMWPGjI8OUwkpjLEn1bB7HUMiwLr24zimlLz3WSRLUjBREcmMVPlq0TTL5cJ7P/RDDDFncQ4dO++cKaSYh67vhzHG5J1zCGyajDM3yW+GoS8J44rQ1CYv6MkQ2KBkGkTnvPeek7oSn65mIlGymjnnHFNIGRCYWcQQgdkBgIgCgE2+H84AMuTCNRcFNCICq3N8zEZoRUtbyJ3iuczOSUrvM+THB5OtyTQCEFQBDQBLgpu7KmBVyXejUydWdGKBb4naB+cr/+L5R3Ze4FyPfCxqZzzx7Snx6M9xt/p3JMtmZ+c8+nIcq1yqff8gxyj3W4H0OQ993LVsovv07xlTjHcqgRPbPfFLcLtqMFloGJz9BceUjHdap/DTJ9XzyQtk2uNkxmFlMSSEcdPWqosYMnCuatOcmQjAQhyBABwZU+G8nzx90iwWaqIqRFRXNQCIGdc192xmKcaUMyGN42gAzjsm1CRdP4xjyPLxPKBv2YFssB3kr3/5xX/9x5s/Xltr7dNnl89/+Mmrl28Ou0M47KUbcBjgyUW7Wvzg3/zw1RdfpHFAyeHQj/24fvqJ91XTgKqOcfzi88+ruqqb1tdN1SyvX3922O6ePnv+yR99Wrcr2u+g2xMBA8T+cH1z0x26Qzf0If3kRz++XLcmOQ6HsetSiG3bLBdXm9XSDPpXL7++vgnZ1pvL588/aRZNHLa7m9/ttm/iGBHdsxefbp682O37w3avaq2nEat/+ufX/8dPf/bz377qQv4mnua7UUt3jmpFh5+z5KymWUFUUkrFVP3YR3G5t5z30nUxpZxSjLHv+77vvfP15RURV02jgCHGMYwp5ZT0yy++4vbKuB6H0QxEBIDewj4/WD/5Nizr+zTEN3PQCKdHqzyfpTwTkxqaOuecd0STwtAAvPdVU7HzohZy7iJ03eHlqzevrg/bQxiNk6EYITrk28UZLAE1hMYUs3YpDZKD5iA5mSWwdOodvm1DzJjxB48/YA764TjoW+07XRQzN029WW/quhERtQxQMv3hcRhiAAZaRh6nRXqAQiirkhExQOlpHv9JVTmNQI6NqSVIqsQnFYHCIzsetQEAjMXkuYyUSrQUECEyMbNn8oiOyTF7Qu9dVTkuBh2OmLByXNVVyRmBoI6JHakKETrPzhF7Z67yy8v9MB4A1CVLMyUyY8aMGd8H5t52xowZMz469rRbLVcYfOv9ouYUgqaMCK6qVM05l3IKKYhKyimG4Nh55533Jd1fTinFICmjOnQCOQKgiRFb1Tj2zESkCpJYwQiNwTN4BkJABTS8zUR3hHfcVJW2OZsBu2axAIA4hEnWIlocV0OboExQjgI8lUkbO3kpEJlBVqGjxFTVih8GM7FjlWIaiMWXo+wiopoS5DyEeKzRu2Z99shWA6AS3Xn0qHgwo1G9t99RtftOod4Uff5QAX13MnZnF4SjucS9He4cxc6meHeKHt/f2f3sK3uMgD7mADylmMTT3wBwNou+q4eC28yBR4fmO0z8FDNbaOY7Z7RpI5xvOePm7OxrmhKl4RlzfV4LNCtEmSBgTGPbNCvEGONuu1dTiVFVNptNVlEw51zTNG0dUgwC4Igc85Orq5iyc0xMRbCdUmqbxoFp312sN9svP08pGREuWl9XRPTYjPdD4c6xk+pnrw9/95tXP3rSXi19/OLL5WZ1efWsaRbbV9cS0n5308W+2WyW6/Xlk2f76zfDYacqjt1uu60Xy7pu6voyhHHsOzUbxzHl3DTtYrGIIQx99+rl79g5A/OVB7Ddfj+8+qrrelX09eKTp390+exFHrsYIpi2TcMEQETODSmnEF6+fi3Im8snT54+M7Nhv43jTQ49akbAP/r0B+uLixiG7fXr/jA8f/5ckb783dd/8fe/+cdff3l9GD5Q7sFvblMkqpuaSVUTAEgWFTWDqmkaV11fX8ecniyuvPNff/31crFo27bPwTm+uLjY7W+YCQFyTsM2NIvVarWq69o7N6o474nIN83l5eX1y89zzk3TtovGOX5njb7dlb//Lfdehz4u4iiUJFtTvAKeLFrNSuw5gIlayiYA/Zhv9odujIdu3O67fRfGKIJoyMeMpwgIhmSAhphAk2oIuc+5SymoJpOsKgB6/P/4HL+7qjNmzPhQePcTdT+i6pGtZgDgvauqSlRUlZkJsMQjATHcDRebhAplAHIcRMiUvZCg5E2+P5I5VuCeXNvMJss0NCiZqB/kPDweDcEI0SMVmbMHrpkbJppcONB755kqpKoooInqylWVd4yOyTlmRu/Ye+ZCQJt5R8xkIEToHLMjZFb26AgInWLuK2nCO1t4xowZM2Z8GMwE9IwZM2Z8dCSXfgW/+nfL/+rZs6vKe01BYkoxElERk6QcY46iElOKY3BExe0OASRnxy6Oo+ZUe48EqnkShCCyr5G9ZpEYJAyiHM2P2K6XdVORQyUDFcMilj0CwbzjRVshCDI1S1tvLsxst91VziFgSqlMM05xmSV5oKnmLCKipkX9WthmMXMlBhJAj9bBZQaSUoKSHwymRDLFvtZSymMYphq9ixF+jH0u0KMBxBQ2+kiRB5+hAeDblLB2rMs9jvk0CTuxrw9oWDvf43b6dY95/SZMZDKc/CuOWYBuvZWPKuXHr/dUo1tTDrs9yAOaHqeSeDaNnNjnBymJ7jHSgCcFtp12u63cI1WC2yrZMbVR8eAmT4QKqIpKDoEdMiWRnMCSWTZH7uLigpEgRiAgJO+cKjhfkfMKkEWrqnbMoIaiU8ZLYFTDGOvF0lX+owV83z+uGgxJ/vGzV3/y6dUPnm1e1Oq4h1VaNC08ebLfHXa7PQyDgoFIXdeby6uqabquizHk0CuIWa6atm0aIjwcDkN/QAQwXS6WbdOkGLr9lp1brpeAFFMaxnGMydftYrlerC6qdhljGvoxp1x5x85DTF3XGxI7FyWZ9+v11eXVs7puDq9fp6ELYR9TRKyunlxU9SKMY9d1OfbL9Yrr9uXr3d//6ov/5+9+/fV1H/M7+OcPxjuW2x0AiQgmzwlCh865qq6c4yQSQ0BE573zHh0DmPeeic2AiBbtIqVgqmaWUnbMiJhTDiGUXst7v1wuV6ulL1JqIkSkbzAKx7On+20Xex4c8e200o+UvrMKND1tAiBWOOgSU3Jc0QGrPDlGMwsxjUkF882u/+rl9fW+G1IGcgYM3pESlHSmxw7WAIVYiAbJXcq7YewlB1CBKWDkfleGx5iTt1zi/XiLGTNm/F54Hw76EfYZ8RSzBN5V3vuh71NKVVWVpHymgMRYhM0wuZOZqYHe/lIDqBllAURiAgBVJZrMNe7Usixg48lNHkxNRaaoJxMFEDVTe8BBIxgW+XNFXDFXTA3hwnHjHCMwgSP0viigqRRwBHXlqykDITlHzEiEZEoGOPkJAU+jH2NQEi2ZLnIIMUd1TbjsFmHuqmbMmDHj+8BMQM+YMWPGR0dYuD+RHyNi3VQ1OWsqA1ORIj8DA1VRlSn7mwLmSKpICFlMRJ5cpRhSGEFFNYvk4mchWQHVNOWcTBMS1HXduOXSr148f/Ls6vLz3XYUVGLRfL9KIfR9j4jeORU77HYp5RSjeo+AsZDjzDYJ5CDFOGXky1lUiYiZmaikPldTxIqIjpnrVESZnfPuxH0zMxGdkqQTvcVk+Vvgnrz5wfwBH8hzTvOwU5H7FslHOfWD87wrw9YjXMujk5l7Vh4PT3OiaG9THZ4f/IxHnkTaBncPeXseu6Wry7mOxznf5XgCnMThJ9IbziaHb1GCn5h/wHurBI+Kr8+XQOwovgZCYKQYxjAMqhkZkIGQDXEYgwGBMRjhcRatMSohADjnQxRTAFEAYGJHJeckIpGIMDsmRwYQo005MD8IA33PkAHPXtxCwT57c/iHz978yadXL368Bgn9brdYQdMuwPkEGMc+x9TrXlJcX175drFwjoa+216b5hRHRKya1lc10gBgKhpDWK82TdMEgr6LYDkMg5glEQNcrS/a5aqqawMahiGFCJKZHJFPYn2I/Rh9VVWNc46WddOuVsQ09t3h+k2Oo2jiyi/Xm/X6coghhD7n1LTN6uJqP8gvP3/117/44h9/87vDmORd8/QPECR+atyTeQtRUeoBM5dsgcMwxGyiSsyAxN43q1UYhhJkXZa72PkQxvKCkkBZACNi5sp77yvvPRGpWlX5qqpVdRzGlNLZhTx6Ofjghd3dag/2fPiIPrbrwzPdX8kxOwqQy/NJSJXjhWeiYm/EyB6YYspdNx768RBSN6Z+SKOYoiOuAE4BMWjToVARE1jIqU+5y6mXPKpGsHyio+5W9467PJ7X7tjVlC7ozrLcjBkzvm/g0ZqrPJ3sHJPr+j7G6L1HYkRC5CmdBsBJDVAyCtrZyMDMMubihwFQMn8YF8flM5QRYCGmS0kEKFS2mWZJ2cxE1eRRsxMDQEAmrrhqKteaNkw1oy8ZCAmcm7IOFgKaixv+8RwiamYEhmBMxQMagMmUEYCYwBi5SLARAVURjT/N+72vPt63MGPGjBkzTpgJ6BkzZsz46HgOLw4buNjGOETCAJ6BTFUYCRBVFcGK+AQRwTMCgQIRKZihgafKoVRU1MaSs0iWIkQ2UAPHZOLIDKlG15hv1st22dZMNE0/zqjIgpjSMIzO+WQQsvTDmFIy0ZwVAEII7Jxz7uRhoWVcbyZZ1IyZvXPEHGPMksUsKzCzqeaccxZTY6dONOekaoSZiIgIiRBRRGLKjyVChwf05d1Xd0ucM6iPan8e+/AOXWhm70xOd49DeQeX8qFpljt89y19fMs+29vovlPG+9sCd5nge94aZzvexurebWM8f3O+6zH2/z2u5/woRESIBkaIzByHYYyxaOZLrL9qVhP2DiuPkcX00HXramkIhlN2RhGTmDQmYlf7KqeklSOmSQGFiIAGqET9fp9j+kDf0Fvb/V6hwyg/++z1j59v/t1Pnm9Auv0+xbS8sHZ98eTpVX/wY9/nlPrhkEXq5aJpF+3lJaqCmajGmLJa0y4q73G5MhEVHccREdm5drEghDfbXcrZ+Wq1WT95+pRdte+6m912GOOyXS3btqk8InZjHLNUTbNeb1brVZIYcs457G6GNAz9YQumddusLy4vLq9U7LA/jCk0q8XVk6dE7c9/+9nf/fKzv//N119dD+nj2Wg/1oaqCgaOmYBUlIicc8M4wv6A7F3libjk7mTv5XAIIZTQcjMbQkiideWJHIQUYlyuVovV8uLyotvbarl0zoUQusNBxVQt5TgMQ4zx9/OAtSMz+0g/9siNc29N6u5uDzWNdjTBSCIxZ3BMSIQEaIBoxNFojNb3absbtvtDN8akYMiCNJlsAAFQMXw3AwHLZkl1VBly7lIeJI8mAigACrdLXidm6k7G04lzRgSwyT8Xj13UFKDy2NrgjP+/4eFv8ccKSPnPE9/YGr/3M4SASN5XzlfhZhtCyFnIFfa2JAUpnfsxy/AphSBMiSSmVA5qagqIkylXsQQ6q6GpqinqlHOwhFghIpScxift87k3153LNDgujqHipMuefvhLD2hWkiCCKgABGZiCkoEZFZkzERCic8SEROCYPRMiuZLN1jF6r74O1doHSIpdvFpX179vC8+YMWPGjPfATEDPmDFjxkeHjvl577q+d0FbDERgoCmH2tdMnHNGRCaCItAjBDRCdI5VtWiKi5akbipAL1lK5DUigoIpSPnAbAyShIDQI/LEDd6buEwfppz7MRBJEOlijklUBFSjmJkNw1BVla80FZ5bFAnNLOdsCghITMWUI8aURRSsCtk5z0zjOKaYHDNgBABVLdOWEgsPAMVAUGKK+dEchPeJm/u2EXcL3b7HB5OZt/Gzdze/JemQ3S387kO9/6ZzPufR2Rc+duqHbTJFyR4ly2dFj6kEz10WT3kTj4KmEx4oxB+9a956ofbOcvc0wneAhISoatHy8uJysd5cv3p5s9vlmEvqueVq6SpGNFUxs6qqlstFvblg0NwfvvryK1/XiEh1bVWd9ruu75hJRBgAAUMYk9HC1C+XKX+VRT5cdqlHv5p73xEqwFc3+7/59Rd//ydP/8efrNaV1xiuf/cF77bL9eXzF58kyS+//t32zSsTsdTD2K42Vz/68U92h77r+mHox6EnxLrylfc55ZTSmzdvnKPlcrler6uq8mNAdk3TtO0ijkM3vN4eDqpwcXl1eXHVOi8pHYa+T+ny+Seb9YVjzqHPfS8pDMMQYgZDv6hSTO3lul4tdt1u3HdhTOIqbC+Xz36w//rl51++/Idffv6Lz17F+57qj7bMe/JK7/1dGCCceFNIKS6W69Vq6ao2hIBIMabDbitA3ns17fveAFzT7Pf7yjvnnKr1fZ9SQqS6quu62d1osddPmoahf/nqJaNcPXu+XC3run7XgtR3uTT7hiY5ez7ebe1RJNGFgx5T6ofharlUtRSTrwmIlNw+aN/Hm123P/R9H8SMnPdVg6pmlrNS8fInp4YZNJgOOfUxDpKC5mgWQROoAcHZd4kwUdZ4220ePwdEICI8Gf1MnQxOJrFi8mi7zPjXgvd8YP7TM87/mScY/C6VL7/3ZV2ImHxV+brKWccxdH3nq9r5yrFllSIIsKOxj6oWxhgRjj4bJz+w8wrblIziNjTKyqGKAwciEaIjUjVRkZxUxVSOfPdjF2hgqjnGoMqOEQEIFTGjFQW0VzRPopCFasdmbFCMnYmYvUPvyFdUe++9Y0ZmcsiOiJmdc955ripYrDtotp2IhJSr/+V//3+/Q/POmDFjxoxvi5mAnjFjxoyPDn+AG+m95ZRTw9KHEFOIMbR165yLYURCPnmPlsF8ya9HdBz6l3hGNDARBQREZGY0ALViqKdqXReyIFGb4sCMhiWZ+X0+EQ1AQUVzGseUxyQimkVyzpNEGTGLSFDVyQpYkhQqGZGAEBHLpmM11AwKUQgARelsUGpVGGhjZiY0NUAslggfGHZ0NP2e8DZt9Xfb99sd5DSRfoTxPf05Y7XOWFI7d6K4F0Rvj0T9vw2P+g98Q61Pr0T0eBsDAOSYVERE0cBXlSccusPNfh9zrpnIOzXdbrery2d1FnZYte2nn36y3e2RERlFpR96X1XEKJJV8zj0Tbtw5Bwi9f161da1/72Jxfe/zOlGHKL+y8vD//l3//xi+Sf/3b+5XLbVMAz9fhejdDEuN5vnLz5ZVG7oDiYpp7jbXgcBdHVV1cToGEE1F00uUtM0KcVhGACQvY9ZlstVSklEDrtdSokdP7u4XG42VdOGkPb7fQrBEFerVVs3aeyHFCXHnJOKEsKyqau6VUNCqlo/hv7N6zc5SN2u1hebuq5fvXz9i5//+qc/+83PPnv1Zv8+Hpnv38TffP8QADMxoeQkY5+TsPNjjFdM3jnJeb+9Tikw03K5XG42u+3W1Jx3lXfM/OTJkxwDAKhmkdg0NaJ1/WF7s40xmhk7t/Tt1eWVd+7502fri8uvDjcfvvt4nyY5SYbfVXwKZDEwBQhJ+jEPlTbEzpGKhSFLH/dd7Po4BkkZjOvJSQkYAA0UEBQJiIAoqA1Z+hi6HDtJ2SSbCZhMPxi3K1UT21Syih7BAHT0j2dEJir9/En/rUVLiQBmqo+wTTNmzPgeUCy1kJCIicjMxjCGEFRUtTyboqanrA9ldHeSQQMA6J0wpynh8rTSrXDy1EIAwFPa4Wk5G1QAxCYLDjMx1aO3xyMgmIy3VCQDZDMiREIgNITCiquhGROBEoKKOVbjjCiacyZmdIwugPfOOUYAQmRER8TsvPOEBK62Zuyw3faDsPsG5/8ZM2bMmPHhMBOLEdcNAAAgAElEQVTQM2bMmPHRIXFsbJXrAdlxzSYikJW8IAOgIAGY2CQ+MbXJDLpEL+IUrQhWQhtVzYoNn2NnKioiklXBDIYhqpJ30UDr2pec42b6kOVBMAIjRlakZMBohoIAoIjsvQPCMs0oLtA5lTlGMdJgQlJVVWXnAEHNjoSnVc6Bc5Njr5pQoarNV56JizZGRdEsfeBR/zEh4entd8S5ivNx9e5/IjHfo1f0zVx28Wp+qwPyWYs9lpn+/WvyrWBlEaWI48e+i2NIY8DJPNYAwDsGVcgZzZi58lWKKQ89eo4hjONYOXaewcRiVBURmSIJzGIIMUbzoKYEWvuqCPZ/72q/99UBAoAYvD6Ev/rV1//2R598+uyyvaibFtHnBBiGHhBpjU27BMC+O6SUGC3udlWzqJu69r6pLoauG/o+xoTMi8Vys9nUTS2qIca+7+u6BtCcs+SsBk3ta+9JtdveHPrRjIm4qev1YgFpjMM+jL2a1csVMqshGBC5umpUchpDP3ZJtFpdrK6uFm0jEr96uf3bX3z2lz///F++vgn5e6UQy5obExNTCAHGEYkc1U3bimrf9wBkkhGMmdk5ZgZEM3WOm7apqmocxy7GccxIuNlcVFUlmlMMopmICZmAyrOxqJtl21a+VrGhHz+kSvK97zh80NM8sutRhCgAIUsfU1Ab1SAbZMmSY8r7QxiCmBEiETlyjCW+Ho72HYgCljUPWfsUDzEMEgfIdnSXhiMBfYd9hkmHPjlvADgsqz+AgI7IOycioopEpWBWLdQUqGWcwl/+MAWoM2b8qwciOsfEBAY5JRVlYiZXNA48GTmfwqdQUU8DgmPKhntHhFuSeRI7Tz/gRDTx3kVqcO4nZid9xaOVnIJdEMxUxDSZIiIQAqEgMBplFSEzIzQhVCEVcUKMkBI5QiIgMmLz0/UaGZZsE8zsnEcgdLW1cXTxkHK1qVQfjcabMWPGjBkfHjMBPWPGjBkfHc96vm6/qNuL5dXlsq1oHFvJR7WuIVox2gA92u6pGgARhhCGoe/7ISdRU1AtThaEyGTOWQjDMPQhjGbAzADkXeMqWyzb9cWKmACygRwn/lTiJQkMQb2nq8vLIeb60CmhqKaU8ciE+MqzcyGE4pKcc1a1ktYOAZkKAW3IR8V0zqqiBt4559yUCr1o38xMlZmJUNTAQNViZIuhe6/2e58AVZtYP7tb8q2J/t59untvH06WHo2Vfyjq/EbjyyIzxPu74qOF76FM507OI+8+0Sku/jZ2/rj3Sf98Nkt81wV+WxLp8fKqmnIutwkAqGgYRxEpPi8qMgn8RU0Ugbz3zntU05RyTjHF2jGagGQ087VDQmYmxDQGIsw5IZEhGGGIUUU/UAz42/xgHpH0GsCQ5F9e93/9L29+9OJy4ehJyxeXyyGlwxDHvjfR1XLhSurAEE0txRStN83W1E3d1JVPyaUUNWfTXDeNr1xIcRzGMYym4hwXZ/h2sWjqWiXvtkM3DIq0vnxR1a0nRNV+v439jWj09aJpFiGrRVPNotA61w193x1iilXVbJ6/aNqWNHTb7ZdffPU3v/zy55+9uT68j/z5g2NyERXJjOB9xc4BmahmyZ6dY0JEYgKAMI6qqqaE0ypZzjnGiGB1UzVNFWMgBkSrKi+pMoNxDEYmWQgQDVPKIaZ3SPPet9LftOWxAtOzCZMDjj3a5eFknQoKEDT3OSWkXqEfQ05BJIuaZDBkJkZERDSd5IqKZIgCGsGGnHZjGLIE06g5gyqg3rd+P1b1JGucRI5IZoTgmTwiAzCSZ9fUdUox5UzMBigGoJpNDckhARVn2JmDnjHj+0X5hUVAosmQAhEAfeUXy6WvanaeEPXo0Hy0TCsCgjuLjqekgncPL0ehdDkCMJNzznT6z0wR0RGrmkiOMUiKAse+7BwEgIAKYFpEDQIQBRVAEDIhIzAiozlHKkIIjlEcZSZPRASOkAmJDFEVxTnmQkADUonYQEQkz94v1t63UBEwQo42S6BnzJgx4/vCTEDPmDFjxkfH1Z/+3Z/+xf/wD8+lapt6vaamNRU8miVMWmGVMs0HmPTOqJZziinFMUhxsC16Z1U0QARmTHEYx34chxMBzVxVvt0levJy8MxgZlPWuXtuv0BIla8EkB3bdEAmIgBUkUL7eu/L7KJEbqoaWpmHMELJAqPF1aGpazMQFcLJDxQAABBKChmzoolGNCxshoFzH/A36N2M8Pkn34EAedte7z7a20Lqz5lKxLv88yOv3kpoodmUjfAtlbi/51ShSVN/x3jjXJF0dlX3LvBDckcppaEfTE0kr5dLz36/vZGUJQsBaNYcU+EXVSGFFEJarTdV3ZikqqrW63W/2+aht+WKmkXdtk3TeO9VZAyh9hU79lVVVbWYbbfbEOOHqP97+incQg0OUf7yV1/9+Plq48U9axbrRe1dFuvHNA49gBVPZ11od+gNKOaY+m4cut67i4vLxWJBiCEElTwOHSIaABN574mJmRSAmderFTvux6EbByS+uNw8/aMXZtjvtjfb3djtNcd2US8vLn2z6HZdEgUFABRJw9iHcSTmZbvarDfD0I+H7cuvX//yn7/6m19++XI7pvfVh73PAs+98u/YYGaWJRNz6xZV1Ywxh5Dbdrlom8pXTFyyZGXJaRhiDKoiKcUYskhIERBXq2XbNl+/fA0Az/gJO+d9PUBISXb7g6taYh7HMYwxRx2HcbFYfRyl/LvWlOjsQbPjghueSZLvtasBiEFUPYQokSwGlWRgiITEyATEZqBmoiKqWc0QMmjSPJj2ol3KQbV4bthkvfNI73lqCkRAAEYkokJAN8ye0IE5wMbzuqlHhIhA7Fxdk6u2XTfEmFSD5JKLrCgmYeagZ8z4XmEAUDK4HhnksuJ1ts41Gb1RGaeVMqo0jR1Pi09E97pHAz4tXZc+hIkcs5qpqoqaKQKWCImUIEsSIZBHflFKbZigIm7YV4A1Uc3kER1iCVphRE/omSvvCuPsPXkqBcA78o6ZkByQA++9c0xYLDhK2Asxs2fHzQKXl1uh4eYGGGF2CJoxY8aM7wszAT1jxowZHx2HKl39r/8e/uO/RyRk8lihCoAhEiCCKk4OoAiAhkeOMCUoEwU95pqTXFICFtqXyTSFFMcYR1UDJFUAIMKqi3y52XlmvGPmeQsDVAU1FIWkkKQImqHIY5JqTplFmdkMRI2QDFRVEYAATRGZiCBL0cxoXdfMZBlVVbJM9iEIhASISDCdoDiZIiARIn1XRvhRPOCgp5aEx6iVhx++x8GnudcpFc+dYx8nZnZaSDibqt2KZI8h7Ld2IXgyUDwTM5+CXu/tc3ZCmyoz8dd2/OxM4Qzn9Z2objsjte6qnk83ykM/gHuwsy/uu3yDZkBATJRC8Jqy59q75y9e9N2BmTw7533O2rQte59VY4qAEMfgfMVMvqratj3cXJsqFJIyadcdPOF6va7b9vUX1ynGzWazWDTRTI7WNt+2nndx/hC9L9NqAEnsn39384+f3/zk2frFysFXX1xeXi4XSyS/3e8lxgEsx9A27ZMnV33Mb65fp34vmiHTVnWxWi2Wy6Zp+sN+7A45J+eberGq10szK0lKnXPMHMaQReqmbdbL9eWlyXDY7m6ut1kMiC6e//HFxUVd1eMQ+64TkbZtmrbaXr+KQ28Ai+X6xfMXQ9eHmzeH/fbzL2/+8udf/eKzN4chfpuGe3dYwLd49NQsi2QR3/iKsBi2pJzKEyMi5FhUDt0hhPjk+RPn+KVZSknN2LuUc4xBrUEiUVmtVk3b9n13OOxDGBFh0ba+WWqKbd3EGILFGONkZP9B+qQHi0mP3jEIQFOr3AYn0PkOp6fzuFZlYAIQ1fbjmIwwZwAjJuccISGxIqqZiCaVmHPMWRHENGruRUbVCJDhnHW5s/4EcBs7cuKoHCETeyI0Y4DWuZqQTSvEZeWfLhYDY4jsqmqxWvt2+dXrN9fdoQtjNkE1AgREPQbtzxz0jBnfJxDxSEBblpxzMa3KZoZEcBqDngYcU1QZIJ46A3u4OFds4qYhTDkCISIRKCBaSSCIt/3Ju1BkEIiVc23dNEgNcet9VYxCjgR0xewdV54Z0TF6x47AITjGynHlHTvyFVe1qyrvvWMCR8xMzrFn9s45IvC1NGu9Przc70E8UP5gDT1jxowZM96JmYCeMWPGjI+O3Qb+w3/4n/80d9vXpNsbUEFUInPMTAxqTEQ8SYxVBAmLTDhLFhFAdOycc6ICCMQsqmBKDCjRWSLQbJKzagbEytdNxa5i7wHpJG/Dk9INFSBmGWI6DHE7jK+3PTmHJTegiakWwXXJYF4uYUqJDiditWQrpClqU4WGCAYiomYIk7pZTY4zmslLmspURzWnPEYh9qapuHwAwC1XegdoD1w4jtHq5c2d+dLRbQKIGBC1hKDaKeQTkQhKBGghWu0BmTgRvueUGcIjc69jfUs2Rrilh84qdszJBcXy+Ky+j2BSItuRaTr9OamVb8mxaZvd3X+ilc+JaDtv1aKYPmtls/NgWDt6v2LZ8+0Ca3vw4tsBwQjBew8BTC2nPA4DTLEAxU5W9/v9htghNk2jWVLKqkqEMcSvv/6aEM1QDBTpzZs3KSWRnFKmut5sNho6ydJ1XfPs6ZOnT5umpd9L2YrvfAvvoKQNYMz2s9++/LNPLv7sB1cLtZvr6/UFVM3ycrPuug7MYog5SUjaLFcXm4u29mnsxzAOIZILaqAiY4hJxAxCitJ3y9VKTRGQkLLIbr+r67quKnOMTG/evGLD4dCHKOuLp1dPnrrKxxi2u9doRgDLtvWVTymlnH1db9pl0676rnv18rUavNnFn31+8xc/+2LbJXmXOuwev3z60O5uffj6m28bM8siAETEIlElkiEBolmKSVVFhJi9c0wkKjEFx84vlm3TImBd1bBcmkHXdYiIhPvdbr/fAwCTE5GqrrjyKafVerVcLJ1hXfffYTHl3vf+tvvgkQ+nhR4zQDTUqZuzO4tRU0E8LlSVhACYAQe1w5gAuSryYmJF16cUcxDTrJJMkkgyzWZWDKBNM4Cca6vPKOY7IujSPeKpAHnm8rMCkkl1wa5lrMFqwqtF+4Ori5iXarBcr+vlStlLjCmGlGJCEuSiZ4cPuuQ4Y8aM9wACGBFVde2cU7XDoTt0h3Ec2SkgarFuvw13KLEKaqqFTkZEUzGAEiEHAGfL2nrsPew05LhlrI8CakdUemyRpJJB7ycmmUZOCoTAhg6JDVFNcspCQIgEiqBk6BwakzIwoRGDFmMOUNJsycS0ZDHMJkkSIYJn9o4zUwQDU8eOmhZFx5QzqudkNltwzJgxY8b3hJmAnjFjxoyPjutf/el/U31y018fZO89mETVaJawcKtmzMzMMqUin1xxzVBUzRSJmJmYQkpiilQMOY0RyAQla06mYIAxGVJdN2HYJwmJivmdHYnSMwpEVGOSKBJSHkKsySGCJAFVlekPGHAhpo9QVUAAJCKwrCdrDjO1XKwAoUxXckyFmYazyM3yohQvVDURiZ0pfx9jn8/+P35ERETTmQimF8cpz+lA7ByeWfvhiT+nU76cQg5rsQc80cnEBGAmikSIeJxZnYLIb7nX0+sjB17Y3SNNX850W4NbcdEpprV8bKda3/LBZ7L4WxzvjqPe6BEe9OTgWJiqEyt/ipMtVuNlwlgIXxEVOd57R6/kj8wSIZJ3rmobEDLQlDWGyI5zyoqiolRcJgBsmriqr2tiBlNVzSmTKQAQoiG0i/bATEeyDIFADVRRDQHqui5Owd+5su9X7K0ctBh88ebw95+9+S9++PzpT1YQrvvDvjHzVdM0Td0uUpJ+GLvtdoPomJt26X2leOj7fowxiYCZIflmWUw6ESmEQETMbGApRTOtfOUrb4RD1+37rqbKu/rq2cXmxacN4u7m9W77RnNaX1xUFSNaHIcQgoFrl6v1ei0ib169iqHPVP/zq8Nf/frVr7/ah/z/sfcuPZIkV7rYeZiZu8cjH5XV3WwOeTV35grSVpiFVoLmVwjQUhvtBOgXCLPVf9BOCwHSVhCg3Vyt7gi4mJnLIWfIITlNNrtZ3V3VVZkZEe5udh5amHtEZFX1u6vIK/iHQmZlhIe7ubm7hdl3vvMd+9Ls5K+rBP+WcGBiInYBEUVkq8I9opiigSNi0zQxplJK3w+iwqbjmHG3b5qWCUoex7F0bUdIUrKbN00TMDrAmEtEcUcAEhHgyMzu/rpR6Ivb961xjCnNz6zPvTknhszPcY0o1cFnZn/UQRxGtUTESIRkQGK2K6UvYzYVt+Km4Fqr0M6jbOWAX3uO50x01WUzIgEQAAM2xE0IDUd3J4DLJl02aRO4Qb9er390dXHoh1F03bbIPLq14C1iw1yIBM0ADOZ6uAsDvWDBWwMCABBR27YxJiQSNVVzgOqfdjbJOQWIajkSqBqCebDS47fBKX51fOU0dL70rYBTTWq3o8X0K6lp9bDo9ct7ntq4m7px9ZxDB7eaiGfoXOfOpgrFAQyMyYnc0YEczFxEkAkRPTAFJkJAMHAjItg32o93EotIiMlhKUK4YMGCBW8JCwG9YMGCBW8cP/rRh89+rqM1rMPFJpmUMh6GfldyrS2mgZmZRcTBichETc0dEKmKowFBXQ99P+SxlEIhECK4RQAGl5IDh5jaUgwgxbR5kcOw36NZAAxACg9KazlWnlnrCsTNKh0rRSvZrOqmBgAxEQKq2UzNSG1Tba2IAgARIpCYukNgCjEAYN/3lX2uJDUzA7iZT0rqcy5YX2JIz/Ea9hmqm2GMlZRHpmpMSkR4ZmRaE06ZudLeeHQ3rNw08dGBuraw1jur3GyM7ABSJEz8+6SiJsTK2NYFmZnW0yDiSWc8LbK8UuM40e7Hs8Ej+4xTnurEhR8rNppVUwl7qSLYuUT5QQcdGe6ZqKofNJ+qz1cl+yQwcjNTN5iPZG4uKqWUkrMUMalFIs9ula+6t78lqpM4c82qVTdVdQDmcLzUiNh2HQc21ZKLiDRdxxxcS+3Y6i/pqqx2fXl5lwKiIxE1LR4OolrXnF6kjFlF7ZtZcJxzcWft/gq+9Qs3uOvlFx8//7tfP/nPfvBvfhAbK2Xc37t7SKvUdrGhYnD3/HO/u2vbtutWIbbtGsci5uqqhMgxxaZVVXAn8EO/q/fndCnd1Sw5mGre70E1rZury5vV1Q1169snv3/x2aeaD+t126Uw5HHoh3HMZrC6uN5c3hDDfv/57v5uvVk9ubef/+7Zf/jgs+e96tdQKn/xKy/Jos9fxFc2eAWIxMyB3RwcQ+DqZ09IqUkhJWJGrLymqU6jTSllGMfQaUoNgo3jICJtm+rOYgiBA0ZTMymFgoLDOOScM7WBiN4ONXpMi6i35LGTcXqzlht88LC7H5nquiGaQwEvABExBFb0sZSd5IPk7Cbg1eYJKruEZ0eYDn76jcedItZ+rCNUIGIABggADVMXQheimxL4Tde9u91cd01yveza9y82z0TuxszjIOM4FqGhT64dUyEqiOKuNSUEFg+OBQveFuoMwZ2Ju65LTcMUiJg4hBiZA3Mgohp/hqlSHwBALYYtpXp0ADPXjLdXdw+1EPI0AzqFzc62QUY0NAdHJyAHADd9aRDAo3p6Ho/MAdwDAjARE6Gjm9bpEREQOkAxNTVFD4GNGYCd3ERBnMhrHeJASIhuiughgKsLhuFud2gvxVFCRnmTYdQFCxYsWHCGhYBesGDBgjeOtPn9X/z3/+e//V/+R0e1kBQUXTrGRlVVpIxY9SkxgrupaBFwiMS1ngq4m6loWbftUWArUg6HAwEQ+ADo7qaWh6wmUsBwFdATAWPVsJx0LQCA4MwUmdA1MW7X7cXlGgD35JWlreyMuXddFzgAgqq6W+UmEbES0KUUDoyAlXYlopRiVUyvUqjVz+vrMcZqqjCJb93BYWcy7EFPsuLXcxJT2jbA0XTDHc3AwdCBABEN3dmNqFLRTExECA7qNXcTpx+I1X2DiInj5DExH2Tmxid3Zkf0qd8qew1V4M0cqnqYGc0qAU1QxUSVqFabHEcI6uJs9sHwuU4PAtqswp69Lvy4gvNj6ipMCzw4SoLONUMPLCXwxCU5AgJVpfTs0Hiyr55P0urRVKSUMDKNOBRwE3vo2fFGgAjupiomhWG6qUKsxghNQGJmVXVVZ649zExA6AhICEi55C5GVcvjGDkRIhOoiAC0FxcrkZSSmZacWeSw3+ec3b7RST3Ug80Nf/juF33wNatZA/jk+f1/+NXH/8V/8ujdP7/qYlAtQ39AcU7Nenu5udje73eliOlBxbqujSk0KQF6jVOYIyM6EhIQegjR3UQEAJrUcGAAEBE1ZcTL1fadm8dNu85Df/v06UcffdglfnR9fXl5AYi3dy8Ou705rNbbx49v4ubi9vOnt3f3GMJqffnkNx//7INPP3jyuXxjM+SvZBZfy02/HoRY+eKcM4J2zUrVYozdqoshSCkhBHC8v79b391ev9ttNptDtxpMmybd3NzsdruxhljEbm/vLi+vYmgAcBgHyRpS17Rt162eySfjOKT0TmjbEPevVtn6znjN3k7FZs/7YRIpuz78e7buwYdPpRu4gAm5BtiXPquMJoNKrs7oM/v8mouCD+mhepCZgCbwGhkMRA0zu0eAiLiN8WK1enRxCSJs+qOb64vIQTIXD0W8H2AcsAwcGYiTaQJvCUvgkWggCuBqoHUMXWTQCxa8HdQph0MIvN1siCjnXL81eAIRMdhUueIYrmYEJkBAcyNCJkbEV59ZxGNWxhQ3fzW9okazTBUB3FTd3eyLnn8zyMX2Pg5mDEYAkTAypcAxcGAi8FxwKCUwBiJmjESBMAEZmCEGRERXFWZgBkIIRIGw5BHRQ+SLzfr66lHz+L0PPr8rvfigGL+/Dl+wYMGCBV+KhYBesGDBgjeOH/7Fv/+H//u/SQ1Hju3V1ksDpWHQ6i4gUtwUEVMMYK6lmCo6BMQ65TeRUkopNRmdObCq5DwyICESYoyNqlZpryoyRwrtdm3rLqaIkA3hlZWDG7gSGCNExkgIiDESESGgmSK6qcZAIRAgErlZdQQGBCBCQmYCYnJzE6UQQghNk1RVRKiJAICIIoKIKcVSwOzkDGhqzEiTgvdkFPGa7sPz/yAAmDuogSO6k0/+GUpQddDMTkZEVCXYxFUdPZuATH6IWkQrP3NMDz3qC6v8WFRlsuCoR6hWiZOLyPFEAKaV22xp4WqGRAjg5kcr5yMBPW07u6vOttHzydf81HMSc2513ZH70ZbjnCg7EvhHAfORjZ7Z99MOK6dFAEDugGjgwUxERBUVz/Jo3xgc3FyLaJGGuItBUO7VVPX2+Yuu7YgopTSOI1ehurubjfc77DpmjCG88847t58/Y+Zms8X1lu7vpEhsUkDX+/vd3d04jqu2bbuO22Z786hddd/NheNh6796g5dpRwc4jPLx5/uf/Obpnz3u/vU7XUoBJJvm+xeflyLtav3+++/f3t7f73fW713HJqWuawBB1Uop4zhIHkWFiNuuvby8qIJfrYkITIiQc3bwFBsi7Pd3z599dn+/E9F117zz/vubi0tw29/d5mE08Ng03apl9BeffHx7d29Aq+2j+xF+8quPf/nh0/uD/GEpwkqchJT0YEMZAJmQ3b3v+3EcOcZhGCrbISJ9P6hJkaIiKlqf/XEYEXG1Wu33B3evQ1MpOY/yKMXQNNSklJoYY9O0sW1STMz8dk7twW944MhhcC4Rxi+6nRy8mA0moHCQcZRSTKvFMxwthqqJ/4MYypFmqnuf7KXJp4G9un0QVs8NTu4t0SrGR5vto4vLR1dXOmYo+d2LTeumu+xmpMZmZEqmZIIIEbxB7IiNeM8lkJAjoROiup8N+AsWLHjDqFNDDqvVCgD6vi85m+nRwmxmqevG54ON16Fgcp8/q17hr+z/QSLbKxz0MfA9CyFeIziYwvG1MraoqNQJqhGZUx2dmMgRDVBsnjQhEAEjGoABGoBN3mWERMS1UGGITCEGIgiRN5fbi0fXq0c3Tw5DyBqTmi8M9IIFCxa8JSwE9IIFCxa8cSDC3/yvfxYI1qvu3fd/iCpQetTihEAIWMW36iWDKjggEajpMJqIlZKH0ZEd2V0QOXAChxBss9kGZg7hwk3NzWptQgTnQpsd3F8/WnV3B8rjrDaZuEtyqDQMAoBrGYfDfgdIuZSqhzGzoqKiXIqIVOvnyhrjjCN5KkXGYWjbtnI34zgOwxBjqrrgUkpdtYiIuzMTAJhZkaKm8HqF3hd0IxzLsbuagNU1xmxBOHHFcGphXTIREFWifrI+5WrVYY5EhECMambmjBgCM7NNOuFJgTzZZOBUa7DWkT9SPHWbSbQ8uXB4/YjPmeyTwTTMG8HMD+PEJJ9kz5PyeeKbcf596oX5g2f08/GzAD7LkY789nwH1mt21FvXd+tJmaMD1nAGEMFk3/HwkK+9IF/27leAiVKMgWh/t4cmMXEI3DQNMec89n3v7rFpuGkFYMzZHMJmDYgmpeTcHw6BGQBMBaXc3d4iQYqBAUCrHbmLikhhNXafgh3fGP6lf36dz54Oqg7Pd8O//8Xv/vMfPVq14b0td02DIez74f72WZFydf34+tEjRxz29yUXBnC31DbMJFKtNkRVkQQJiHBy3lDJpbRtG2MMITg4Ebr70PfjOCDoep1u3ns3dKnPw9AP989fmHnXdev1umnT089+fziMoenWN+9kan76k1/9/T9/9PHT229FP3/lZ74J8+jVsUdDoC6uV+tNHqVJCRxEavlBBvSuay6vLtdXl58/e4qASGim4zAMw1BKQbCaOR5jjExd2zWp1dITETAjhxA4hCBSoIipqZbvjRudqJwzRudI1LwUEMSXP3cejnN//X1r7tnUsvTuBVzd9QFtfRwtq4bazw+FZ28RICOCOQHUVHVwCIRNoC7wCumyaW426x88evzo8hqKiF8AACAASURBVLJru/3dXd7JCjE5ZIDiRghNaiIxATAiICaClqkLwRETUy0SRoAIfhyHFyxY8FYwubk1basq+/1hGMciAoBE7m4iLjZZcBxHBnc/I6ldJt8LOh9MAADAjttXF7HXpE9V76QJ4mavnTwgAAHUuRoRgxm6M1GMoU2xjTExp0CBKTKFwIGQEQg9MAbmwBACBWZCCIFiDE0KKYUUuWlS28SUUghEjDEyprYfchEDQEhbuu3fSMcvWLBgwYJXsBDQCxYsWPA2QEhYUx4xmBYviu7ogEdu2MkwIle3OvSAlFau6lJCkUbETN0diThwrRPopoSOBJWjcEBXAzUQt/bqPm7fff/d1bOD3Y0Ok33F0W6iiIwlU2AsrGZjLkAs6mI60eEKZtiP4uBmxsxICI5gAG5qOlcWJHAHTllBsxTDnLUoFJMqrKkVwxRNxMyMZDKsZUIkDjGIZP8aRrMwS4zheB7nVblmOmV6veaFOgACOvrMnyP6ZHJaaSF1QiAgO1pfmAGSHSs2IgCgAmC1LXVAAPPqnuGVOT6yy36WUV99VAEAvJY4nPt90iX6OcE027uencLxlP3EQs9mHdMH3e3s07Py+bj2m9aSlc4+7Wfyg4QH3grVcByQiAOpg4t9tffvd7UpmKIEREjk4Goqqn3fP7q6DkREpKJ1EVzrJJZSrAi2DRBaNRwP0dwkl5C0lFyTfEWkjaFbtRzY3c0BYpDSq8ib9hV5iNccywEOWX715PZvP3j2eJsu29W64bZrDFz3/bC/uydaXV5fXm4C+bDfqamMauDMARFSim5Ooubm5ipWk6MNoEhJngChOs+Au4r2Qx9ivH78uF13MTV393f7fV+KguNqvdlsOkI/7G4Pu70aba6uKXVPPrn7m3/4zS8+fPZin7/vzjrysN9Q/eoeQ4yEBKiiZspMzORuDgbg1dsnhNC17R0TEgFiyQUcyL3kbEdmhBAJQwgxBFPPh54xAUDbtgaupnWM/dot+6JHAF9RLM8+OnDMTzh1wrfuZ4fqaOEKptMIj+g4MzkAVqNNx+F/MvWojx0AuHtNtYlMiF5z1cGdANddd7PdPr646BA2MVy17WW3apl06Mv93Xh3J21ksNL3MmZFrkO9FHHzWi2MAAJhZA5EPCVhfKH4ccGCL8D364fz9vHWbvWX4p340osceL3umMmslu6YbZUdzLzW0Dj/vJkROOCcOeZUg+vofpqJIDoQHEPkDs7HUDxYraGNRHWa6G5uUmq8+zXuTnVcIMTI3AQOgSM6EzQhNCE0gRNzYIqMkSkGmgd7i0yROTDGwDEyI8TATZNCoFCp6moGV3KeeHT0WA6+H4bsgPCLe7hJb+aiLFiwYMGCl7EQ0AsWLFjwNuAIiGKZ+vuD9DsbduDKRIRo4EiEhGaOCEyMSMgMMQChMwIwciTz2VkYqbogm7oLgLibEyIzqqAoknkb2027vbpIbatH+mFqCACAqpRaI5zJHIooIKiDuZu7TQ59WEkud2fHKo6uuZQijmiIBKBESMSiBipZ3MzN0bSqih0BiNHFRLzmxZsagLcpYjX2nQU3X6cXT/9FgknUSwAACJOKd5Ycw2yZilR9rSdDjKNsmWZ1sUOlYyrJS44nwCwenJ06Jv8KOnsXj5zy0WLDj6Tw1MZJgXy2ujtZccDsOf0SOzezzpMEqTqV1BOZjnHOYZ0d7kGPIZwTXTgfegbMpo1ujkhIzGxuNpci+3Lt83eCg5ubunWrLoDnIY/DsNvt3C3GJsZg7lJKEqlXyM20P2BKwIE5dl2X+0PNv0XiNjV3DiJFXZCJQy15D0DkMYlqEal16v5AmHpfDD7v9W9//cmfvbf90XXaRA1N6rrG3Xe7/vbFUwG7fnSz3a6JIA+DSBnHzKQxhiY1SGTuWlRVARCZpgGBAxKpq5uhuZuXUkR0e3H56OaxMX3+9OmLF89zLil126ub7cWmbXl3+/zF82eR0nq1jqn5/H7/Dz/7l3/3k1///vND/noxoW/VCedEyZcfZeJSmYNJHg7D0Pe5SAgxpUZMVM0R+mHY73bb67FNTXUYRiRTTSEF5DFLluIhmJlorSBKSKRq4+7AEM396OEOVB3GvylJ/ppzOQ9hwWmMc5iplzkU9J1g7o5ux2F9ijfV0gDHxvmcPOKT6TwiIdVAFEIVOwc0i4RdSgQYOVxdXLx//ej962tSadw2jC0RqhyGUfd72e9h3Dqhi0guGuWUYu+TeBLdGSFUomself9jZxMX/CHwH+9d85bZ54qXOej64DFz0zTgoLXYNVK1dQY3ACfklyyqCNFO+WRTCWcRrRVKfc7TMkBAIHz5oO6gpiLKzExIsxxBpQBUxvp1FQYQmCgypxQapITI5Im54co+YyCKDHEqpIhMANVEjrEqoyMTY90ACRxMXVxNrIC7qZuaKZHFshMYDYEpX2F6lr/Pq7FgwYIFC74YCwG9YMGCBW8FKAVpv+8//t1v874fd7cyHpomxRQdIMTIIYzjWE0qYkwhBGI2MxUxkaryq3X0iEmLqIiZuBezkiU7ODKhGwMEIE1PP7rTIY/2BRyHuZkdXfRAVWeiAt285EJElXEmpKpdAYfIwdEMKYRQmVARUVVVq3YT8/5OcmAkcoBcis3+EhSIiByhOl2AG4DNjM1LxM9RK0cPVqFE1R8bkCqR7OhnzCtO6yY6/kB3MEQmCFW2TXisNnbMPGXmuiqqXDHNrtF4ymWf2kQ4p9a/TECDwxkTM63SHiS8z51zRtbgLIJ+4Lcx09dnXDiAI4I7HndwdspQc+eP/h1nu6r7q2eFblTJ36osPvNs9KMp9puGz/9KKS0juIuIiHZdJyL7/b7vB2biEKhtIQYiWq3X3Wpd1VZx1bWHZnf7fHN93W4voF1dbC8+ceAYm5R07J9+9umYxyZEzRmHITCfW5b8AeEAav6rj5/+00c3f/bOas28Hz57/O67TdOqgR76+9vn7n55eXl5ebEPUcacc64XCgljiF1KUqQ/HMQkcjA3AGiaJqXkpmLm6iamZhcXl5vNVou8ePrik0+exJRuHt1cXj1qV2sONPR343AgIk7p6tFNL/bb3z75+1/85p9++2Q35DdG1X8DRqbe4mZm6ipuWkqWwCmGJoZIjjFG1cmlVEX6Q59LqcbvZpAC1zKGDrDPOaUUmGJMzNG0RyKOXGXyd3d361Vq2m42iv92p/byx8510MeBzM9e+V5wkjfDHLU6Uc9z5Iuq1WsljhzAUQ0REIjBG6J1jKDSxfjO9aN116271dXm4rLrNjHuPn+WD7t7GT2lJsYGQ8cMMbUxNYyQ0jiMYmYIIaYmtcxsU7DOAJwIcVJNTsn1+EoO/4IFC94QkIiYEJ2ZESGXPIyDipgpEQHUCh8Tv3z+wQfTC0RCdATmY33k6V2CY2B7msUgERPVP4mcqLLXNkXo61j4uoLABBARUwoxJY4R1AwxMiMxIDmgOSoYOdR/WPP+ANQcQdxpyrhDyATDyIQ1xa1+GszMEZGDxwSut4esbQSLSP5Xf/1v39gVWLBgwYIFD7AQ0AsWLFjwNhBHoQYJCAFjihqDZiJm5jBJQfPYDwdRrRswkRtMhnoTV+w1Z5KIxmEoOZsqERC5qFT9r0oBNQYsDHf3rmNBc5ocGB4yuxP5W71/K9tKROwAimbigTEEAgQiIiYTAwAGA4KqXDb3WiwRnPionZmkvASRa1E/IgJAN/NT9vcsUVaR1IzDqCI2GUp8kfLwpfTSmVmZyV2kE8VCU2nDWS9OhDUn3IwJA02v1YqFMBPQhFg9rM2NiZEQTgXh5wPCzBjPPPKJ6/VzGbTNiuRJKTS5Rx/bfvrtXqXa52V8zghodwckqK4hs6v1LLUGgDP2+NgWB0AgIJhU16eqh5OQqVoL12pgZjr7NrqZVz766AbyhUzRkVv7ljwSIpipiKSm6e9vu8hd111eXR7290S8Wa3d4X4Y6hUJxIF5P+wdydxlGPf3Lz784F8utxsdx/7Z09gOVkZzV/UiGlXJITA3TdM0qYZaZr7/7eOccpzowf2o//Avn/zwqnl08SfvNHbY95vtxfbiilP7/O75i9un5nJ9fbPdbna2c8fqnw4Oh/3u9rYAABKOw9h1bUqJOZRS3B2RxKyIgnrTNCGE3d1tdYJOTKv1ZrXexCZK7p9++tl+fy+qsV3dvPvjUeDjJ0//6Z9/+7N//s3z3VhJ3D88HFQ152yNNYG5aZnjbt/f3d81qyY24cWLF2baNM16ve7abne/iylmFTNrmqZtmq7ttORcSg20NE1i5mpS36S03l50622/3wFACMFUh2EQUf/GZ+8PhqbXvHHa4OEA982E1l+F87DTlO0x1xCbxeTzeIUOhBQCR8Ltqru5uGiINm37ztWjFEIkbkJszPzQy35vh30AhVp/FRHV0MzVAKnmxJhqyVlKERXwqVYYETNUBTQSITnisQjt93ziCxYs+AK4u1mIIYaYYhqGcRyz2ZzMVacIQK95Gufw/RSofxhKh3nagXhOVE8/juWWp+/dI0NtDuazCc/Lx8Q5wcwRxE1NxVyMIlshTkxMwAYExgyRiScPaGCCwBgIGJEJCZ0RmRFpyiGsrmyqBsScGgLmiGrgxmiFePV9d/qCBQsWLPhCLAT0ggULFrwN3Pyrfxp/+uf9uxeb9ZoQc+KxTSmlGIO6lZKHPCAjGDiYmqhCGQVm7UmtEMdEVZTsbipiZkwxhsAhArq7juripdTs9OLkwAABQCY97WnG7wamXsUvgScqPHIAABEBZWYKgSZFdooaVNXclBCZOEY2MwFDQyKKMcK00tHaZk4RHMwMq9moHfW8x3ULkjUy5j7EkjO4fRGJc2wyADzYxv1UZQuQmWa18rlyebawADBUwqmKzqyApuk9cERkYgcnoBAYz+sK1g1gYrx9Yp8dAXyysLAqajZzd1NTmE5xWpBVrfTswnHmtTHvajqdl5P46y8Dr4bT81azhfOJHT6Xf9diXzQR8UeH6GMm7cyeK1a5tlmlkMzMVI+aaHh9iuzLzfvWqKtCV0MAMGCmOBOpMJtV53EEpDIM5s7EZRw8JSSMTWpSY2qmCoQQOe9GDoGZkTmsVo9ubvq7Z2qmACEl0bu5xtIfFhMRqQYffnb70w+f//kPH1/+MB0OvaivLy6urq7aVffks0/7wwDwYtWtQ4gJkJlVtZRSVMyMCJnDZrOpoRwHM7daQdQBmDmkuGo7lTIOh5LHQIFiWG82IYXDYdffvSi5LznHtru8vsHQvHhx/5tP737+4bNffvRsFHudOu2745tHLLAGlrCIkOUYoUhBQhEZ80gBAzEBqlrO4zgOxOTmplqjWQjY932tZtk0jRTZ7w55zEwUQlBVyVlidvPNdkvEHELTNBz4W2X8fxEHfawKCnh6gs+F0d8ZZ+7+AFBlgSf2mYAQGbCWMmREAkd3JI8xNE3TxnBzuf3xu++sU3vRdZertZVShlFzVhEtRfY7LGOInAADQBEBVVfTIgJcRw83E5E8jnkcbW3EjMy1WiszBWYmwlrJdqk/uGDBW4S7u2poU5NS0zR+ezeO2R9SyYhThP78g8fZU90J2BR9Pwt51/2f5gl4fK2auVl1dEMzmoLz/uo85yWguYlKNnUxUAPwxJMHdGBiArOC6DEgEzIigweiwBgJAiETEgATxkBEQARMyFxj3k4INRPDqLpeY9P8UA4vvpeuXrBgwYIFXwcLAb1gwYIFbwPr9dMf/w//1z/+H/9TWq2bENeJbdMBgLtlkdjExrv1dosI1fjCDbRInedP6mKfks2Z+S41/eGgZtVFumhWUwdODTJFY2u7S2nj++/j5Ud3jJ+8auhaiuaigUPXhfV6o2oARMxuVgnl2fWh1m4pdSFi5grVLxhtKkWI5pZzRsLq8Ve9O3Baa5gWRZwEcW42jrkSoe5eSqmrlFn+fFae78vh7ipQ2dVae8tMbZZfz+Tz5N08+zu7GU0k0MnVgggQcXbLgElhTjT5XUzmqfVAXjnu2tKXmlMV5T6T1jPvPe+LTn+ectD93I7Z5mXcyRBj6hOYWwzT22d2qz6/gSfMMnM4vXDcyVR/DGuJISKczFjU3ax6qahOLXr9MvGcRvz2MsZa2j4GVimrlAKiFBn6PjCHEERkHEcAMFFXdVMAiCkiMwAQUoqpW60sj6bqZoRIXE9r6prazz4z1Ignx5U/Bjj47aH8+sndz373/M/e/VGLo8oOEFbr9cXlZZ/l9vb+sB9K1q7tEIGIOJAYMkTmQIgxhtVqlfOoZl5EVQOHkAIGBAAmcjcpqurMsVtvUtc1TaOlHO5v+7tbBEgprdfbtmkPh8Onz+9/9sGn//DBp5/eDW/E/LmeNMBXBZleBiISB1cvpahaKQpAiOjmUqRtGgAvOU9xCwcpUmvolZxHwFKKqlLgNrWIPI45j5kQQwhmPg4DcwOI280WAYm4Sam6tXyf543zY31yynjJjeP7OxQiAxIiVWHgKX4JbsaITYjkXgma7WZ9dXGxatLjy4s/efcxDCMXgbu70h/GYQCFJsQmBIgB0LrAq7aJMUlfOIS2bZsmEVgp2RFDim3XhSbhOKibqmTVXLJCHflrnKQy468xWlqwYMEbRYypbduUUi5ld7+TXESkOlJMBmt1yDjDlK3jNUo9qQZCYDjFxo/lRE+zBa/1DInq1E7FakLWMTvstU/+8cDmlscRc1EEtBr+dwsBPTAmpnCcDp+DEBgpIE3FCREDYwgYmEKkFDkGDpGbpmnarm1XFqJx8/vPnx0c4ZPPwo9+9D108YIFCxYs+HpYCOgFCxYseBt49F/+v7/5f/47TIlCiE2LpNwGc1d3NnWoZcEdiTgErBSjqld21WHySjarjAzHsBrWrpWHdJ33YKpmbgbcXrYjv9+ni4uPj2v+82W/u6uaiDohIRatLDDV19W82ndCXVuITPYUZm6GMKmDVRUm4bOd1M1qpGYO5i4qlQVm4kDm7jlXWTe5e8mTt/U3FsVV4wo4mljUFx/QonXBUzeaXZH9gXDHEdHNKr98JH0dEafzOjK2J8MNIzx15JGn8plKhlncPfHNswv1xH7OCkg7LsWOnLVNBPZrRJLoD5xd/chyTx0A56xeVYXXXFec+enT4WCuA+ZmJqUii4hKZZ/N/FV/xrlHX34FvjWVFAI3KaUYwQ0JmakMNgzDql01KZmqFAEDohBTiikFZnGgGIkQa7gCgZnNTIbBmyHFoCpKaCKy39/d3ppIQLIi2vezd80fCQHtAFAcnrzY/+SDT//i37x/dROil3HY73d3GGPbrkTgsOtLlpxvQ6Bq8cyBkbhexJq0UI1tqn0KEVXrHlXVUoaxEFCMDccQV6t2vTaXPPQ6jgHYADarizathv1wdzf+7pPnf//Lj3722097eaPM4Ev9/5WHOqr2j4OPO1oIIYQIiCGGeRTCpm13u30NGtUajIE5ptRIUjdETimJGyHB9PBXZyNjJiJ2nyJQ3/yMvhGxfmRqvuduJpgqlTISExIiuxPgVAAQwAEC0iqmSJSY2pSuLy6uLi8C2GWTtoRDyXoY1EyHwXIm5IDYxDCYuirHiZcvKuYOhDX+Z2YwmW5wjeaZO7ipmUgx5Mlzv15HsFoL8WHXLViw4HvEuUHWlHnWdd1qtSImVc0ln2Lkk1+PH+cnVbYMMHmzncLr4HjSQhyV0F6fepiF0V49zeaZ1jHuO80O54SsV3EcDhiJkQiASKtIIAVMgRJjIgyEQMwEMVAMHAgDYmJKzIk5Bk6BmCAETJFDoBg5JY6BU4pt1zZNG1Ijjhrbu10qWf0v/yv49NM3dzEWLFiwYMFLWAjoBQsWLHgbQIS/+9//VQg2qqSA0QghMDMzp2rMiRN5CURQBOxYPhABAExBBdSACGJM6w5UQbUUUVVOkZmIKt3KQAGoeXavT8a43W5tph3xjEVEBDc77A/OVHLu+9EcQ3QAV7Uxj0QUmJHIzUSUg1WxjKmCeTCrVDVMqxGrstMqXzUzYlEzVSUmAgTPtRb6TLiqu0uRXNT85Aj6DZhorATwrP6tJNVxTTXZXZzpoasYsLqgPpAL1+N6deE4GkPXJdaskqbjbmvXnewxZri7O58ftFquTpLkyn0iuFXfiOrtPbtFO7i7mk08fj3I6Urhg7/n0z8qo+Fk6wEwV1CcWwX1kpmazv7OXtXOpjax/3aUYYMfqe1ZrjkbT5/0m5Orx1GR/W2IJJy8X0IT07Pff3R9sd1uLgLz73772zLmzXp9cXFxf+hTStS0TbtKIb548eL200+vbm5i12QZc84BPGJU0/3+YJKLaNs0MQZmRgcZMxCXvh+fPh0OKGfWIn9QnNpwfxh+9fGzv/+XT95bv3vTUtfEbpU+ffIxYFqtL9fvbG5vb4v0OWd3VxVVI4opJkDMJY/Ph8PhEAITcYwJEUsuvUgpI6gGYqe06lZp1e7Gfvf0s1WbAmPXrT00q/Wm6Vb3h/7Jp88KdD//zZN//t2zZ3fjHwH7fC6xd3cbc4aATbsKHPrDAYibtllfbEPbfPbJ7xEJAJEopNS0zXq1enE4HA6Hy0fvXFxduY4qQ39/v7/v//Rf/+n68sKk3N/d5lIQseakl2F48eLF9dU2AojKMAz+zSxIvop6Phsk7JWXvhdUq5KJdyZkRHIgAAJLHANRQATzxLxpmlUTN017ud5cX1xs16vd3echD7qj8cVz2feO5KpszgEDeAAv/UFLbgOLqDocxmEoGcyKSgDDGukzq3VoZ8kkIIKoKp0KDxIxYq03S0dqbOGgFyz4XvFqdAcRcbPZbDdbdHQzgFqQkGsyDQCY+/HrvZRSRKFWxaj08bHwICIxuzvolCeFiIEZCacZzVmQHxHr/BYAECEQyZyn8iVAxLZpViFGADBhsMTURG44NESRKRIycQzcxJBiSDE0zJEpEiXmFCgGJrQYqW1DDBSYYuIQOASOMQKSqYA7pQRm0yzm3Xe/32uwYMGCBQu+BAsBvWDBggVvCYexeJ/Hkre39zDuUs2cdyOu7s4EE1tKJoLgKcRZeTtRiQRuZkUkMAdi4loZvJaqAyRIKQKQiBePz3vo+71ZYYRXq2pVkz5VZeYQAuBYGWQHQEfiQETADABAyJFCjLXeFMx0JQKEdORbyVwBgImTu5mLObsDQiAGADefHZkJANAdEXPJiDgMA5RyEv1+HUaiOmtUm4UTnzx137l54TnXTBM16zOffFI7VmftKoV2N4eZN6Ez8hppNtGeHDl8djQ9kySfncPEzNjslXFserX2qBwyT/Lnmf6u18ammo1HUTfizPhODto0d/x8pPobABBpcoCdG4MIzJOxNSKoSCnFRjNzFXWwuWpitf+YXUoeUGdTU74vCfHsM+KIuL3Yutl+tytZdrtdm5LkvNsfRAQAMOfD3e1uv1uv1xeXl4iYh4HMHt88fvbpJ26euq69vNLDvm0bMxvHzB1c39zcP/29i6Zu1bz3g6e6qyvhPyqIwfPd+O9++i//6fsXqz9ZrQDubl9E5n44jETp4vq99955cftid39fpJSiKSUiNtNxGHIe27YNIQCAu9V7UkSkFC1KgAoQEolL3t/d7e6LyHhI2+12vd5Y4+3ldR7Hw1D6jJ/cD3/7j7/5+LPn36T23reIOpwIka+32YNXqml7fS72+116HlPb7HY7c+tWbUqx3++Hfuj7Qc3aLq3Wq0N/2O/3pZT6IPSHg2sSEVMtZRiGQ85jyOMwDtUXqHofvan75ES9fN/sMwIhRqJQzU+xEtBO6AFplWIbUuJADpu2ee/RdUIIbsFhbbpSGceR0TiGNQdv2wg45jEXYfCAkJibGIopuhNWKyWs46QUQQJidiR1LyJFREwxMKfkZm3THEWVMNkfvRxHW7BgwRvAOQ3tAJhSbNqGA5tZKQLzDKdO+ciMAgNiLdoRYjC1SkBPu7O5hgSzuzHRsTgGEta5y6xudpyj+GfNMZvr6D5MGXkwGCYK6xjb2LSBgwM5MXkTOAVqAiXiSBiImhgCMaHX9I5AjOBmZgi1JASgF1fVjOiEjuiTIRmRuYsDpxZWw24YHBsA+OlPf/rmrsSCBQsWLHgJCwG9YMGCBW8JQy7iMEhfxsJ536KMw1BKBnSs1VWqlg1RVRCgidHN3WwmWQHBTaWUEohDCBSCA6qjmQEYoMcUwHAcS8H2XsJ+J1oyzf4b53AHM1DTSNg0TTgMDlYZbQdkC8dVRM2YjjERkc/FZUSkUkJQ9YdEZlVhOmmRXSofTZW2rgIZhGlJgwD1s5qEOSCxm8Kkpvt63NZRjjypu19+58Q+w1kxwqk811H9PLPCRMSMiGbminiukgacl00nn8MZVv86ej8/6ODKT5ub25SofiyPSDQ3Es+y8udPTjQ/nPrB5yTXk+kHwnExN+XDHrlqPxLQMz89nw4hITozmRETKRqCm897OPl54DnDeNY6n++l78ii6ey9knMmdwAQkWHsQ+Cua5koMLddR8RQq+qFoGohMBK6o7tXk2h3NxHLBQBijGBmpmYGbjw9UO4lm8orLiJ/eDjAYZRffvTipx++ePe626yCHQ6BIyIPwz4X6VYbcI8pVWrgqMonmu6gwAHARUSkEBMzEXMAYEQkUpPcF3UFsMDs9T7iwEiHfjjs9odBDoX/7pe/++VHz28P+W2JUb/+hUBAjDGCeynZxMw9cKglWMFTiilwiDGGyO4mKqcMBoCu7Z67l1IAYb1e1+BE3w+llJSSmampm4FDShERSykll++5AmM91zcsvUeAgBgR0T0SRUJCY+BEdNW1227dpQ5Etk364eUlavZxtGFcmaxd91IQPIoFYoxA7iZkgIQYJlFhBBWu3vFIdQz3UEdDRGJAmrM4aqhgGvRDCGowceJE7EZTYxfV84IFbxQvjbEeY4wxmnkuknM2MwQ6d9KY/2MIyMQvP6M4x5/nmQICIZ6yp04bHudWD1tj86ZfFeKuzAAAIABJREFU0mgmSiFOpYTdmSAQhBBCjXsRAYEjAQXAWqvQ3NzVEYzAM2FgDFMqoAEoIiA6odUZnYOLuYC3m0uGdBiLNOl//qu/+su//Mvv1NkLFixYsOCbYCGgFyxYsOAtQczJXQhj07QJNsGHJg5DX0o2mHz3ANEAq2uClKJFbGZymdFUEYwIhlxUHYnGLFkkcAB0AFGzkmUYCneXhTd3B8j9gU7Ovyc4gIGLGoewaZr9YYAizOyAAKhmVRLs7pVfDiEQkVWf4MqLG04SGPSZTnRzY2IknLwg0FXFzMzUzQHQA7s5uAUO5kaTOy9OZtLoX5eeMDeyypNW11egE9WDgAYO7nUtRERo6FVHiVPmJVbfQwAAUHEVQSI4inrcRRXq+eGsD561OxOhfEZFf+HKarK8sIkvnxnzyiDOBDlOFLJPZs80sep0/ADNsuTZD7r+fNCAc012/YnHRpr75O8yibpjE5GACKUUEznWgaxGLbO66XQeL90/eHrt29BJZiYqauZMIiXFCIgihQhDYEZi5hgjMgEShxhjEu1NLXAgJhMspdTuc1XNuZTxuOYm9HHs1Qq6u2bL/ZgHna7mHxfE/Nk+/92vn/z4vc2jzdV1BI7YNE0pduj7/b7frDdImGIC8HEcFSSl2LapaxMSMwd36/s+5+zgTdsiYslFSkakLDlLBoCmaWNqmq5rmhbAx/4w9IOI9wWf3I1/848f/P7FfpBvxLx+Rw7Rv8bNM2UexMCetZSCgWKINVGAm6bZbFbrFSGMeRjzsGaMMc4pCy4i3dV14FDv5K5rQ4iBANDVtBpqH+uNxhARoIx5HAazbyIE/+rTfPN0q4MjsDs7gFnDsYuB3YJDF+L7lxePLx9dbi76uzs27UwtjzIeWErnaUN+D+COCdhrZEcLOTAhE0XiyJxCQI0pBAZ0MxCNzKFpUowMbkZ1BI4xxaaJOddgZCnFVOu41aTUNrLvB5wMU+ZMkgULFrxxuDvEyEx4OPSHfd/3YxElYvdaohnc3FQcXFUJCWkqg0Fnps8AgIihVhd0Q6SpmsUcQT+mnL22CQB+dJeecrfOqndU1GoZ7q6mpI7gzmQC4uAOgkYIjJYVAiKCu0mtUczoTECT3hnAJ8Y5Bk6RU+IUAzOZgzo4MYdGIWQ2Qvhv/+u/+N/++q/fZP8vWLBgwYIHWAjoBQsWLHhLQERFCCE8fnyzQm28l7ISLVpL+x1d9hBVREVNpOSipQBAYObAUjKYEc31uAD7fhxzjjECurmWXEqRbuXcbpVXvKJHl92qBS0g5/6jk5mDi4iqMnHO4zgWRDbAyn3XynnV5o9mZraUXFcciGhWZSYTB0pEDm6qhoaI6lbPxdTcHQnBK9NKqmKq1XdCVb2uFghOKt6vhBuAg6GjA/JEJwvM5hNHg2KAc/0vVuXwg/I7p82nV86E0bWGXxUVz7uCWkVrFgxN2501G4/C4+NibHr/wbnhQ8B8QDj6Kz9UYePJU2PauZ9Zf/jMMU9ZrrNSezq6uaGZmcNUnBAAAAzdj5GJB4opP/vPwy559f1vBwdXM3VP61V/a4DIHIgolzyOAxMVyaruiA5exfWBg5qROzkgYmpS7g8AXms9jjkXKQyA6BzQQVULOgAaMUgpJ4b9jwkOIA4/++CTP/3B9kc37dX7TbNeNU3bAlMYPn/67LCHEONmvYkx1oQJQm+bddt1CI4czVzN+nFwgNQ0zOwAw9ADqKgBEDOH2GwvLrY3j0Dt7umzF589lWLt5nqX/R8//OzvfvnhXZ/fbu/g2X9evYmObjWIAMRoLoyeUnKnw3gI7rFt0nYbQ1SVu7vb+/vd4x9Q03Ui4m5MrKrqFjgE4rFkkRJj7Nq436f6/MYQU4xMDAhmCuZObu6vhOq+Kd42t1rHIQZoEDnGq67bdk2D2DGvY3p8eXHRtQ1hP/RWcogEKmyqWhJoS5gAxQ3UaklBlUkV7tXCX0RFpJTs3jSNE5dS1AEAcymRERANQG0Kl6pKHYRU1VSdAN1PCSpz3dQ/rkyEBQv+/46UUghhHEcRwZkshuMXO04TiDrTs2q4MRUhBICpAMRpbKwpWXN22JF6pqmS4Vwa96wBU42L10bq5y8BU5VxzObgIKoRUYmkUC1wQlNZDW9CCESIQOAEztVlAx2JiCmEKQpJiMwUAjETMDkRuDMRpRiaFgKRBHf88TuP3ly3L1iwYMGCV7EQ0AsWLFjwluDojCElurjcXgT33hDaOlOu2YnVooGQtEKk5Cy5EtAUmHIupoLuxISAbtAPw5hLiAzopppzETU14rRSbi8Kvff41xdr6u8M9MzAof50L1LMLBKZm1pdIoCpmSiQo1P1BEQHAzH3POaqog2BAUArD+5m7gFDJVKr3rdqhBXA1JAwYhUnnpwBj74T05pl8qL42vSN22SlTOg+eY1Wq5J5RXQ0Gj6r4+dW9c8nXrc2gCZ/6sryuhkAEtNM/QIcTZtn/hfRAQjPCzvCTBUf+WwihNMqD452HacTP24M8ICAnjnnWdKJL4vYsXLQZ+zz7BFSOehZKQ1ewxX1+rq5gVXJk7v5g4r1037RcdZifylR9B3lnUhEhFByjHEcRiJpuzaGWKQoQBFxIFArOedhKCUX0bDZuGrOg+Ssomo6lhLGkZrV5eX17WefiImqaSk5j4F53a1X681+HFITmfmPk/ZygBf7/PMPn//5D69//O6f8FiIQxu5a+N2u97vey+WS5gd3kW1PH/+uT+HwCGEGFOj4MScc/79k4+rPhgBVBUQmTk1zXqzvri4sCLPn3/++Wef2Vi6bour7ZMnT//2nz54etdn/eORpL50l6MBMnPCxMy3t/fIqPr/sfcuS5IcWZbYfamauXtEZCYyARSmumcow2khZ9Ei/AWK8BvmI7jkniItwh2/gBtuuO0PmP0IR4RkS4+wq6ofVV1d1Y16NIBEviLC3cxU74MLNXP3yEwACSCRBTTtAEhkuJuZq6mZW6gePfccm273VWQYBjO/vLzc7XYAWGtt+mViFpHr58/VlEViGp98/vmHH3yolcdxQsRSJohwNdMKYGa11npxdfXwwXs5p6Xg/BvgD9ONAZGIdin1Kb9/efngYrtB3DBvJd3fbLMImPlhH2WSiw26YRi6pogEKG2hLbw9ft0MIgjA3Rv73AhojDA1YDQ1DUAgVW3BhwDo7rXWqtVUw71xPRCBEQTQnrqnNT84PZ2+P7fdihV/IHx3KzLRCtGYqOs6kdQI6OOa/J3tFv+cJm6gFpt8DIRoq3bNaefoZT8XwM11aHQa72BghJ9Sr9sieBuHvP4hiRABbqYW1RwAyCyQHMkFm+VU8w8jBEzmTASQhEQ4J2lmHUkoZ8lJmkX0HPVBKDQfAQBIhPuu220qEBVz5HhNQsqKFStWrPgOsRLQK1asWPHOgAal1lTGcRKrN9c5JZHkMMtHWASRAYmEMaEwJlXQCmZtMp9ydnM3bUYKANBtt76Y97mZuZuDA5H0If29SB8+un91kT8/FKgOzTh4mXe4xzRNxHz//v33h+GwH4lSqarVcksNJ6qqTJxzJkKP6PtuEbdEo2Br8xOkZhlNiLnRoQChalZrIBFzzovY0Dz1uWlaAEBVh/FQplH1S+ZgMTttnMfXEAIQIAHNPhVAd2hlmE1LZzeJo3oY53eOpPPMgNPC+MKp4JSa5S4znblfzJOlE228tOikqT6B4K5D9UkadCbRPr177qV49s6JA3/pfpp3x1gKWlvE4VEuPbtqL1mIbZ3DzaxqKR4ebr5Yv5zfGkvI4aJY/MLr8s2xsOruiCBJ3OL2dh8RXdclZnfYFwUIERYRIiZ0OxwCAdwjfByHWspuu93du58u7988fuJBXdp0/Y7Sxv261tj7KNsx33+QkiOgv/nyxtc/nW/TGxbw8WfPf/ZPT/7kX3/g42CHw+Vuu91cPnr0cLMZbm5upmmIMCJKzLW6q7l7sNVpslqAONQCQjVyzoxoaoTIIinnlJO5PX/+/DAOh8PgyN3l9uq9D3//Qn/+T5/84jef1O+yX74Yx+/AUYL/8gbhrqYtvWoqkykys7m6WyM0u67bXWxFuFnM55Q2m41NY6211mrM7o4AzNJ3iITDMJRpYuYup5SEGGn+goKZllKqVkJ6pSVfcgrfCyBgl/P9i93Di4sfv//wwa6P4eDDROMkkjMxEmUMx0gcVitoFWAwsKoIQQzEQEEQ1NyBmMDVoFn/IBFLEmkK6LZyJCml1AljuDMLi8x2QABqxogiknNSJCEKd3dviWF0/iA+c9WfyzICv+x5c37GX73ZGxbUvONDvfnRvp949931hniTD3334vu3+Ilf9+6ae0OY+77b9Btmfn59fRgOU6lI4uBucx2XexATIpqeliLNTKu2iA8Rbu5r8EovN2LX3Nv4K5rhG6GZw2Lx0dhlCJtr1wAAfP76I5wfEwHCPQCaRTVQiMjsCMTUdBgJQxCYsOskJxbCLO1dzElyl5JQEsrCSMjMXZe7rutyTomJOIii3zwbpmeTTWDgb/7AX7FixYoVbwErAb1ixYoV7wphCFJqefr540lsev5JlzpJ2WefZU4pE3FjRgHRCcANwwkCAxDA3N3MzZmpkYyEjEusHyAxExCEzdylMHaZN1mE6sttAfDwqZRSJlVtlA0zNccMgNn4wM0a1a1qEd7ktB4GTSoLcXQ2cLNwbzOQhQSdHYeZeY5TX5jrxkO0gD6Ao8EEngX9vdpeONJ8iIREs3SZFuKZF8fkNumZC0LhqHNeVNALTU2ACIRAeLK7uOvdgR6OCLNNNZ4ok4jj3Ol1RPLLguUltmc+6knuvBTQz1sdJdtx5I5fNu549aezqtiF1Qs4OgnMpDISAiBDAKIrQgRVAsCjkQie/4fH3c6MGl9/Rb4pTsbZpOp913PmcRjMrJYqPUtK4oDE0O44N2YiDANEkcR9yrkwIzFJkq7rNlsiYWImBgd0RKTwUFWKqLWq2ZcnIH0LfFuKIQCe3U5//9unP/nV44f/7YNtKRMNAJw9ui6NI09TqbV0XSs+JmExN2wFE8xm7t5sTHj2akdnZkmJiVT1MBxy7qZaiKi/2KVuU9P257/9h7/6xW8+eXr7dlP3vuZ5v9p1pxeXegBgopRyls4dxhLMzMIIqKpEHBFaq6pqrWamqsyKRBe7i/2Tx4fDodTS7y63220hnIbMRNZiGxFSSokFW9AltwcVfT+V8l8GBGHZdd0Hu+17XdohTqp1mqIapozMJEkAgHmTkpqiqoMzMxEj4dGKBwEigIgAyQOIGvMzpw8udRZzpUoEmIWpulsrbW9e/O1XFUKYuUG4OwQQUWZmVSwwP2DOL/33vce/1fLS///wB+mu9QK9FkFMfdflLiPhoaUFhCNEM0tuAw0iZCJcsigQAFviNCHhnG0LgIhtsHenYooYAQDV20DMPRoBHQ6BMR/W3XyRUL98BAAABCCAzLKRlAETUkJkhMzUJ2FGIRSmxJyFBCExZqZGNItQFp45aOGUiDBEqBNuLUmMgsAQHAGuZoBd52bECIWCVwJ6xYoVK94pVgJ6xYoVK94RQp15Gid9/PizG6zT889ySkmyewA0AjpxU4khRrhaheZkJyzMRNRqzCNippkiZHmPmZmFCM1jrAZkIIqiEJoTMb6s60MAd5+m6XA43NzcPHv2fBimTX9xshRelLMpZUSaptHNWaRadTdiakpnnHUvaKpzfhciwTyfaezzHCxzZAANArS9UmttcTeIGEhziedrgbEwpYGExALYPooAm0rnXAJ9pn2mVo9JR8EyLqJhBKDF5OJkdNHKSM9YYkRo9FTES90TZyKe46Qq7m4xs7wnM4+T9m8hnGcq+vx/y4HudgguUuvlIiIuJiJLPez5BnEkdhyi3UutTpYYgeDoNDBXxp88Ne5aaC8ipVPtLd5hzr8J5pLbWWKOwMKp7zbc+EStWmvT0QOQe6gqMlJOVhUQkLgFY0ZEHUcex65PiOBhqhWnwawSwjHc0efb7/tbbDtV/93jm7/6xe//u//q0YOu94BxHMdp6vq+6zMzlVJVK+dOkhARu3Rdl3Iy99vbvdrYbfrtxQ4RtdSAYGZEVNOqVc02m22HXQBISpL63z09/OXPf/OzX//z7fSS+8YX6ZHfLr78+PO7p28yERExC4DP56V1GIdxHKdpTNB5OESM41inqtVELDz6vheWdjxmSZKkhyFnAAj3Mk3mRkSSBJsWesnnhFMUKt5t1feUKEVAJOpEHuS0caOh+u3ehwHNofSQEiARgDBvcjYAChiHkUUkZ0QEb88abE83ImpptO2XEeH85FRTt2bZ425m5hE+lamUyiLUVgQB2tJoeNRSKqBUBcSUUi9JSgWcAB0gcPXfWLHiuwczdV3KKQHAcDio6vHB2qoZcAlEvruaflzWp/mBIMvS+120UjYTa0OsY4grokIEMyGSm5kdNRBxepaeOHBggD6li82uA8xImYkJE1PH3AychSgxZaYs1CXOOWEYE+QkOXEWTswsSBRuSghETePgpZRa64AoiBYxRYjGtRph8j75oXzHV2DFihUrVtzBSkCvWLFixTtCTXvb930vV7v06OpR2WZhYU5uPk6llJJSImYERsJwB6U2AZDUhI14GKZaC4sIErEQACB6RJirB1YDBPco1YMcxTlDEr642DFPAPpSe8J9HIZxHNUKQhC+TK8gNN898Nnew9FnW+Q2zTgyoU0c50veVACYW7PlmINnFu0zs0SE1doIjFjklz6r694I4W5Qm+8GIAMCEKE3LnmmoU9nQeiLP0ib9sxcNAYC2EzftlnQSQt9rgmOCEQlopMk+U7KzpmHxtwZrR79ZLCMZzM6WMTjMB982eNscnesTL3TJ8tptXYSEsxmIGcbxVnjzuydA2IWhwO6qZY6jWMt1c2OOtOjC8dRkX0mRQU4cZOtEXH28temkhrl7w7msNlcuOowjBBwsdtdXl6WaTwcDpNFlIpdh8weUafiIl4rTCVcD4cDYUTYuL+uqjmn8OoAtY6GXuvoVpAQ0VPK3YaRyL8rre9bOGwAvNiPP//N45///ubDq0cXHaOXaTrsD7cfffTjzWZ7c3N9c3NLjBSsVSPg6v693HelVj/sq9er7YP7D98bh2GcRguLCFWtWgPi8urq/v37wzTe3Oz3t4cNbv/ml7/76S9/+7sn16+YP7+tLjq/K76Etz2yuq+9ixo/AmExjlMtIZwAoZRyfXNbLVT95ub2Akk4pZzdHRGYyD0Ow2EahpTTvXv3xmnSwOEwZkb0APd+07t7KUW1tPUMtRjHaRxGM58rIV6j0vuewiOeH4bnia0T5stMNHhk5pxy32VCHKepTiUwtGqZpvEwjGPRnbabRNXCwiPUzMyROBAjwtxVq5kiQs6ZmZt/vojknFNOYEp15qckJRFpy43MJMFdzghIKeWuy8QVEJmRqDlK/bCNKFas+IEgSbq8vOxybkt0ZkZMxNS45VPt19lwrkFEckrnC+pf63NlfhSwmZr63d8GZ+wzAAAQYibapHzRbbpAQRBCRhDGxEQYhMAIbfQZEOoOWs0UIlIpLNQKpBa3aEhMmyxzPRlqG7gJU7AocdxMBw8VnJ4bb1cmZMWKFSveKdbH7ooVK1a8Iyhq+dEnH9z8uEtysbkoWloRtKk1r82UErEgEBJGOBtjABGysAgDQs6ZiFJKfd+JiDeJKJ4bQ2CEEwIQElNOfHmxffjgfkrXANN5YxAAIqZp0qpEtN1uiBNTMpv9go+Wx40DmuuwCYkEAJY886AlKb0pjk8q34DG+sIyg2nbpCQBoWYBQBHBbaKC4EddzFcTmhEB5oBwrPeGcPRmAz2zy3PzEdHBl0CaNs9aCOj5YI2JXlL/mpxwoaoRAcDDj/rlRVt8/APOpm6zsenRSeOcfT52+3IcOlcRx3FWdtxtefWOXOiMJ6e7oY53eicA3I/HOarC28HmzLVa1TT8ZPx8Mv+IxR4kzs72Dr4tGdfWNiSJbDY6Ps+IATiMwzgOzI8udhe1WhxGiBj3B51KzrnnDseRIlAkLNrFyjkR435/czigMGamnNP2vftCPl0/8RZ9RhTx8urL9xDV4vPr8T//1a9+/N5u011eCjFzrfXp0ydJkvu8RFRrqdUA8Pr2utM+AAGRUwr3aZxKqS3vaRwPgQiIueu73O0P+9v93iw4724r/OTvf/OPv396GOt3yQHi6db9Gtuf/YzEzG4uLP3FZUqbWvXm9lqS3H/0wXsf/shqbcQoRoB73/W73S5KdUA3G8bhxYsX++trFrm89+D6xfW2E0Tc9Btzy5IwQmudpmkq5f7V5XZ30W8Uif4gltjfBhFxW8rNOOlUUJ0ZUY0CEpEQBgD4XIQBgODQSgrUDCDmJ0OAL0mmbfWqFQ2Y2eIc7ziHjLXfM0iL/REgBIQ351bEJoUOQI8wRENo5q+BBIRAtHh4fH8J/RUr/sUgiex2OxGZyz7MEYiIifisKmseNRxVCB5BAMTs7hGuasfx00tPR1wWz9suJ576uOIes/nGawZ2y5o3AgqyIHE7oIdZBEYYghBhIARhKCEzVYKWMdhKmhiBuTmBOAAQAkEwYWZq/kGA0J5hOSXuNrTZarVDAHawuYLh+gcwNlixYsWKf0lYCegVK1aseEcoF7cPb98TCK9mZm4AYY5uqgTR5ZxyZuKjeTFABx6zWR9BID64d78J0FJKiFhrbSTAcdAfgWpeqiIK567f7n706OFHH7zf508A9i+1JyJK0QDo+/69h+9Nk9YSpdRaLcKbnA2gVTE6dhgtUV2ImNy92a5Kkjm2q01rmJuzM7YgdUR3bwJqVSWiruuQyCPMrRHTdZrG4QDRKEUM9K/gn+/ohANo3j4QwCnA51RBBGLCaNFzs8sHwBJ+h4g422u0xh8JasTTBSCiJipvZh1L6Sq9VKB/Hj7YrC0gZheP5WjzZmdm06erACdiGs9O7+Vy1+Uz5w0J6a5hwh25crg3z25shDoiIbXaeTcNCHM7rTScOva4nhGvfPJrrsQb04t3NeIAHu7hEaZlP+1fpO1FSomQaq37/b45F0vKeHlF+/1UpsPh8N7D90jEx8lNwZWZtXopJXPKuY+A2/pCgKza7bPr4TCG4XZ70ffbw2G/v51KKX4n/PEtsoxvx7YiAIaif/3rT372b3/8/r3N9pEkStldtbYYqGGs0xBd16c+uXuZxmmcEHGqRafp9uaFmQIARHS5dzNiliQ5dwAwjdM0TZI3CvLTX/z2Jz//+PPnt+bfuOVfed1fa2Hx6r4vHefOjxFeVZHZ3IdxqDWEU3uq1GG4efLEVHPOLZFymiYWns2dORHi9fV1i0gFNVXd7rbmOgzDOAymNk0lIiSlnJKbjdOIw2EaJ/MfHh8RAJP5YF4C3QLCQw3CgtBUmVMWybkTROEEKZeUPPYeEYg5d6iGzGgKEIAYsJS8sLdKFzcfx2m7uxDmiDDVMhXvMgESUQSoWilFrS6JuFFND+M0IcWFHabpUFRzH6en3IoVK747xFFpnIS3/YaQzFxVzRxidteBeYzRFpgCAKAN+QDMjJqD1RxarMJMzPEFibXmThFB1HJfEcF9lim4GXjgK7stC+KAAATARG4+DZOao1m4ATgT5MTYPJHQGYEJhYkICSKl1ITPwsSMABHu4epa3RTMck4piTC3lfSU0vYKLnZXGmjhGxJg+1//43/8zq7CihUrVqx4DVYCesWKFSveEf7Df/jz//N/+x8ppgPo0ycw3TyncCKECDPz8L7vc+okyX5/W6syc5eyMJda9of9YThst7u+7xvnYqa11oBgoq7rRDKLREA1n0pFpCTZpgPpdG/b9dJExtFY1OMkAhHDQ9Xc3M1b+TkzaXWr6i0SHWfLiGhGukAYNIuaEdwcCFjY3VXV1BYdMJhZi0RvG8/MUa24uIU2MItIan69GHFmXPwFOFbHn6gMnPMEZw3zHScNXIhjmEnk5R1aRNLgiDS7jQBAE30vnxUQhPOOzceC6MRhL6YdZ3ofXAwmjj13bOzZpgBwR0K90NPHFxZRO9wx4sC7W83HPzHr82bRZOzu7hCx5Ek251Ydx7GU4qdQvjge7hVu6Euo5+PGb0JfvmL0EGBmpUxWJgBHmpWRbZKMIs0cIBYf7JnH7zqfCiCwiIgUM1XtKW22l+M4hQNL7tKmREyTmkMEITH1PWLB04T32+BL5Plfrdz/SqjF59fDT3/96b/58PKjh+/fu9j1Xffs2TOtJfFm03cURIAEgIhq7k0Jbg7uWkuZUtd1KaVopvIiKSVC3N/uh3FEQgf+5Nnh//7Zr371+ye3w/StbXhfuzue/RmvvPJNPqGtYxWbIEOLCQw3qMXMmJlFmIWITGvMayygVftN33WdjkOpdRiHH330I3Cdhr25HQ6H+w8vmKUVoktzKkUS4STpm7TzD40AmCw+L/VHAfeoJQmQEBNimJvPIsYyzV98j1Ct0zSN42gRXWwAaTbfgLa+hcycUkopQVgWQSSLtpDVTLkRwpvZSwAGoDlW90ENATQQcg7ECmgsIBBMQAxEgRhv48uyYsWKL0YAACF2XX///n1mHg6H29vbthBba20EdCtxgMXGi8jaOMKsqYmp6RvcXAPQfC50OP4DYGoA4O7zcKctY89xC1gRw8zN2hgEjkOO5bcBETbveTOdouw1kgeFQ/isenYlgkaYM4IABqA4AKGqhRsjghkwULPsyCltcmbOSVKiJJxSkiRJJKfcXd7vHzz87PbweL9PQ63dSoOsWLFixbvG+uRdsWLFincHrGiMMOmt7XW/J3QhYgJVczcCRzeIdLh5MY4jMV9sdznl/X7/7PmzF9cv7t+/v93uck5qqlpLKQDBLNvtrus3krJ5NAU0AAhTGfc67nshOZo1NIY0lqxzRDMr46hqptZK+93DW+U1hM9V1U0LE+7uQWAnVw0PbzJhbSGEsah0du/ZAAAgAElEQVSJPZr8hRb3i7aLqiLRQuhCLAXdc6vuuA1/ST8iAgEB4EzHwXLMhRE+uiQ3043ZGXpWAiNBE1vPkWOxJPEsBz+qkWc18Gzh0bptORodNdW4KI2PDDOcaOZYrC2W4J8z1nw5l/mcZx552SjiFKMHx31OTTt5cpx92vzpROQex253c21ur1arqltLJfxCl16ENwkJ++bKXwRw81I0giV17q5WEKDFabaMTbPJD/swlSQ5J1MNgHZHSRIEMHcEyrnr+10p5gbhwClvUt7f7vcOpVT16He7nMd2l75VvHr635ZWC4Di8IuPP/2bj+791z++ev9qJ4lExGp1s12/gcBpnGqtxMyAm20fATCOwsQsKaVNvyGicRxFpDn5VIvxMJnZZre9Hv0XHz/+i7/7+PPrsbxi//yd4WsZcdxB409ZCEXcyM0hHAiScL/pAQKRmKSVa7SMVrP5xK4urm7LtH/xvNbCZl3OBDL2vUgahuGDLguzqWnVLCmllHPKOYnwK2b439XZvV0Mbp+M078z544SMwEl4cSsAKYKEe0r04ogWl180zbOGYQQjuARfCSYWsorNAcmdgcDnx9jrbDdXbV6RABqgAZMFoeqGFA9TJIhWERFVCQNMIDGPv/gTE5WrPjh4HzAgCmly8sLRJymaX84VK0QoGaIgQCqGh6wlHy5e/Mwa/VpBiYijZ5ulPRpiNYGKcvvwLPFbITwNnIEhEZOg7m7LcuJcdxwXq9vo0AzdS0IEcAQhAsr7h6IAMgIQASIRMxEiQkxmEAIE0NiFMEucZ9Tn2XTdRe7DRMwY3u2dznl1KXtRbp3f4i4KeUmJyoVVqxYsWLFu8VKQK9YsWLFu4NNvZDjbsopdxcXHWNOTIRmqmo8ZzjhdrdpNhfEHIgOkLt8dXXFLKrVrBITABAhoJCIAU5qNYqaq7sbRPhU/DAOt/tStTZqmGCmI8Nnqgzd6zTtb/fEYua1llrdW2V+U59ic/fz2d8ZCdwC3Myae0Pj9WKcyWMmbhQHRCvA9EYmImJjqOdjAhzdIUy1TBO4H5W4eGcK9RogEZHMhC5xI35jSR888tDM3OxBFusMPIYRHuXC1Ayf22GX/ecfF2Z3eXfebFYAHWdfbSYWjeE5hgIiztrnM0V3RLSefeUcj9vgGfsVcIwojGZ3eHaG86cu/PTJs/vYxIhoztpIyLMgElUxPGCpjW2rBNB8SuBcIvyG7PPxVL4WZnILKUl/YeOL4TBwQEq83Ww2XYdEnGQDYGXMklPiCK+lxP4magnmcKtVAYJFWBIQE/FUyosXpbu4uP+j9y4v7j/95HdVNcximiJcTdsU+tvhVbbxpdN/Cxz07z+//sk//P7ffLB5uP1oC8Plpo+cdapalQBqGc0j5Y6ZHz16pKrx9OlYxs2m3243/Sabmpl1XVd1qtURpe82Xc4K8Nmnz376D//8d7/5fF/1a7bytYsN513xqufGm2zwZYiAJt4NjyzCKZeih6kkSMSc+g4JEElVm/k1Iu73+2kqu4ur+/fu3bu8vP3808P+dhjH++9/ZO61lgjouo6ZtBYzLaXsb2/bOo2Z1lKmacIvbOVXnuMfEoeqH9/c3r5fmbd932F4Eum7rgTuq6WcM3OX86GOaopMqev67UZyKqrqpuFVq5q2pQt316rTNI3TqGWCcJZkROEexBHg7s1B2z0sYpjKZDZ53EwlzGvAwWFCdPO92r5WVZtqVXM/PtRWEfSKFW8ZARDLYjm4eyAws7mVMk1lcg8kWYYuyMzA8xgoIrQqLtGv7u7mbWhBjOEBgLMt27I0fyKgm/Y52rq8LMv9AIAYblrrMMSr605xtBxDBGz1KAzAGNjMnQlTQiIgQiZMwlm4T6kTTkzCJIyJcdPJJktKJExCBGFZeNNlAAew8KqTep0KjZ3HpttM08FMvZpB944uy4oVK1asWLAS0CtWrFjxDlHTNPUXV8+73e7exSMBFQrEMFVTJeHG5+bdTms1c+ZExJuri1qrqUaT/jbyEwlFPMADkAWQolXlR0BghINbWPXeHmreXW1yx4fiACcSqQ3+S63DcLi4vIqIm5u9SCIks2YRPLPCiM2CAyKCGAPDzKDpZpgBwFp9JYATzXKYAA+PxkUHIaK5zj6DMVdgBsBcHx6BROEOiyXxV9B4MyGLAWcG2D5nIJ4roJ0cADAQCQjAPQB8dsdodCti4DEkZ6aol485jx2c2dmAWax9PETAYhSxKJ1Pmy8/HnXPZ2GFTT8ecKJ+4VTbejzRs/+OjHhrxxyluHhInx14ESPF0tHtR/dwR2iV9Tk8tHlju0W81N6vRQx9AxYpIJAACamOFSyudhcc8ezJ4+sXz+/fv0KiMk2OlB492j9+fNjfEuHl1SWlJOauOg0jIubcjeN4GIbNvUddt93tdr1gJppubl68eJFzv91kQri9vt7v91OzA/5OcLxb3w4X6QAff/L0J7+6/NM/+aP3E/IwXvb95mK3v9k7ESJFaCllu91GRFM+ExMi5pwi4jAMt7c34zRut93FxVWfN7VYqXo7xT99ev23//jp7aDfuie+gez3G3ROtBjJ4wIYBHRdp1ZfPHvm5ughRA5AxF3XC6fcdbXrcs5V9cX1taptNttAevbsWc754b0rQg6PlNIwDtc3N5coDjEMAxJ0u4uuy12Xvnj16/vCNb8Wxf15qc+m6cU0TuOYCJlZ3YvFWIuaCeESKXgkfualrOWJHapmaa6+Z5GcMzMFc9d1khIAckoegIQsAi4iEgyckgKUgALoAK30fgDcm5fDtK86qBWrY6lV1cO/fH1xxYoV3xKICBHMvOm7q6vLUutUilZzc5JAoFiipCEcPIh4Xhfy8Nn+a66dOtLT0fJImo4BFiHzgmijO28lE7BUfYW7h/trvvGzyxhQgCBmThlZEBKiIBKiECTGJMiEzJiE27+dUBLKzMyUhESwz9InEUYREiIAYqLFcY6RWvVeAEY1p6mMpXigjfcyrQroFStWrHjXWAnoFStWrHh3sKnvPthDx9znq0eP0CbwAhCuGmaSEjIBRu/mFu7RSp0RcTb0dQcIInQPEt7sLqtFUXNAC/AI83lUjxDgFlo3k4/p+sHDq/53T7CWmZJctGcRoFXHabr3QNhgmqacck6pNnlseEAQMTMDhLmbWixK41muwgwQAA7As+0gEyG1iYy7zzHkAIIMALPEGWluRgRCVRVkwaiv0ci8Dm1iBLg4IDcOZTG0OJLQAIC++FN4c87wxSoDEJf8vbkENJo/RzPoaGQTHWPfG/Xks2y7tZOQAhotP6vEsbHRCzPdhNFwPO2TohoX95HFduRY2LqIm09c1x1Ha4DA9mlEOHPli+v1UrO6pM57QADSopNe5oyEJCJN+xwR1uwaz7IPv7jjz1nqb6fzjfAAc28e4aoa4d5cxd2ab626QS3h5u5qVsrkqm1SPeu7AUREcobcIY5dzhjq7gkgpeRupRQDzPfu06eTe3xnBDS8XWoyAJ7dlp//5tlf/OKT/+FPP4w4jIeDEhOEamVizFnNx3F8/PhxznmaJlUFiMOwj4BaLXWdiGx2FyxctbhFUPr486c/+/Wnv/7d5zZ7wJ+v8rwkcH6T03mbnPuXfEat1SUiwNxLmVDm0or29ZnGkXOWlETk9uaGiYQJIAix6zIxEVHucre7unfvHjMXG5o1TUp5u9lcXFwkTpvtlgjHaRyG8QtCtn4AsIiD2ZNx+mx/4MN+kxOnlM0mtbFMxZQJq6lHNKvWZsbRbOIBoNkMqZuZeURTR6acmAWSd30nOYUji4Q5ADAzpsQpBRBKqhEFYEQUoECqgPvAm2IHm0aP0WwoZazaGvCGz/kVK1Z8YyBil2W32VxdXT1+8qSUqSkACAlFwsPMEDHC3B2Imgn+cV8CQp6NNojIAwJ8WR9HPB8ytF1oLqs7qyNrzK/5LD14BQGtMi8RbVLukTJEh5QIhTAxSvPWYBKmLJyEhYnJhSFxsIRwJAYCcw9HcqcgJiT3GK0K8+KoFBhB4aE27Q9lUjC8BzD6D9Lxf8WKFSt+0FgJ6BUrVqx4d/jv/+zP/vP//j/VKT5/vif4xKchdEIKZk7Mue8QwbxqreaOQSl1ImnmRmmmPk01pcSSAEk2mYkDsBlbNFLTzQgBCYOgn/xg3fuPHl7sPvvkxQRLouCxSc0xo+/ydrObJu27XjhZoyHciflojhyzPmZWMDMSE7UJjKrmnIlITQlnEbGZqemR7GjEqkd4QOMgmJiYdKrX1y+mMla3xhG+Xv4cdyvjFwlm43yXV3Dh3zEg3HzRHRMiOvhJzrx4QDcOFuAYD7gIqNtmy0cte505b8ybnTTKs8EGNofTo9vzqcS0/XHca9kJjtQwADRn6ZMJSJsHtjCgNrNrDDfYvAiwKMbblG9WLh0pZ1/I8cVtAxFppu2Jmn024syZvztSCAOgqpaqKGIAWmsgiHDOmYU9LMCRGMwgXE21FkRqVDVCCAIRaUSLuQ+tROBu4aqmyY0ZW7Snu0k4zm4lb6HlX7XB2+nESf13n9/8P3/9T//+jx/s7ouElqnklAAhZQmgKFVVb66v+80mIIjIzGIaAxBRtrstAKactdbxMGCkF9V/+qtPf/brTx9fj2e1099AxfxFJ/j2meh2H7vPtzEipJQsKhN3Xb/pNwe+UbXUUU4JAQ+HYZqm2WilPW3c1cw9UkoXu10dR1Wdm4vITMJiYiklIiDitmT0g8bTafpslH/FwsTQlg8JaH5QRy3VA4A4kMyjaC1VHYKTEJFFpJQQsVYdx7ERQ6rVVIdxTIEVsJqqRQQchsGsDqUWh/AYU7o1PwSgmXqMFi/GaV/KaDZZTKqjFjWzJrpcsWLF28ed0gIi2m62Xd9F+DiMZaqbzYY45W6DTG1FFomgqQ0QECmJmJmZHZ8YbWWKmVXV3QBgXky/O0Q6/1Ifo4PdzVytqiK61iVS+ayaLAABhKnLebvd7pg3ABkpMyUiYRQMRBciIRRGbGUaEAYO4BZoCqYUbhDe5ZSSMFOLMIHAlFiYkLyNBQCZNqPxde03wdnitoeLd3RlVqxYsWLFgpWAXrFixYp3CnMwJyvl9gZ03NfxFtxylr7v5TB4aCmDqkaAcCISRI5wJmJuqWJhaimnlHO6voWUgqVZGdNCXhIgCxEhMLqyBDy4vLy62GI8eYlgCQBVnYYh1FKft33XSvwTMzNGzMQEAFgTyiG6u0cQERMzMRKEu6qKSKNEjwQ0M7NxLCzonHITHk2sbc4tTc6BmREJW6Lga/mJE/t8l4MGAHSMY5zNIgeeadmjLzQAgkcc069myhjbcTGgxbZH68A43+wceGTvX07pWzwyjuplXBp70jIvGubj5O3kfHGk05d0xiUGjJCJWm8jERK2RQaHAAy8Y+sxH/NYYu8YgR4R5hEBzVMFmqx7doGGU5e9ESv09pijADNXVWB2j8AgIhEWQWGaqrqb9B0KI6Gbulvfd8zsbuEG1FI1AwDA1MaDe53KkAkRXLWYKUAwE4bZcHDTdnO+tfZ/xwiAF4fxb3/96X/5+08e/elHm90G/WCmKMwiEUhozByIEYGEKSUzRc5ERMwppVorQNSqh6EQ88efXf/kH37/q39+NtYfEP8X7RsJEOEODP1mU0p4eJaUU2oC5yQiLG3hbZpKuBNRRJSp1FrNTM3HYTAPVTWzVgNhZlpVVU1NtXZdFhER+cHcIl+AJ+P0mfBHm9wc8Gl57CbmJAJt3YxofoZR2yTmVwDaiiMREhMSHgmtgAgMD6jm1d0BJnfzqICjm7lngAHwEGBVi8OodjNOg2oNL+pFtZi2YNvX3H9xp+TjzfAmd/EbHvMtfiHe4lP0zasQ3hbe4r3/Fnv+e/uNfPeN/8pPbEvf86CCCbe73Xa7Y5ZhGPf7g3kg4xJtPJfKtSgPXMqv5lEctfCMl0DHsc1SqLUkXZyW1CHCAwMcAGMOLjwlfMQcfrwoqAOAiYWlrYA7gEGoOTi4gWIghFBwG/uEhRuTEzkSMCI3lXY4hCcp8xDJ57FZ36UupxajCBCSGBHdHYAiOMD/lz//87d6gVasWLFixVdjJaBXrFix4t2CnZhUoSrU4sN+9HHfddk3NSBKGQ+HG3cn4r7b1Gq1akQws4jMlCEiETVHCfOwAGRiFuGETJJS33VJmJkiwnkzTHy56a52WwLwM60tAAREmcrh+rYcDkIM1hRyyElmHS0aMRNRKZO7M7OZhQeRuIgzM5G7m1kpxdwBFiMLIgBobzWOLHyWNDZljaoakZuVUmqt4dFo9FZcf6fHlrkNAh1ndIt9RkQ4teLPJg9ulaCLaQU3BSBA42GPfh3HPiAkFnZzM4NGmjPHUpZ+lxbBRmzNdrRHA2gARFpkzkfvDTjfHefo92P96jJHPE+Ph1NY4rxZszBkbgQ0EeHsT90mcRHQ2rl0VxwF0C07yB3APYgiEA3A3cyMANvU0Oxoun06l3cDRGBGJvZqbiod58TTwfb7W9Va61Tq1OUeCLuc+67zMrSllc12A+6mZZpK1Xp9/QLT5r3N5fXNC3fLm77fdMBUywhhxCltNnT/Pv7mNqXUCLh3cHLLX75Vf1aNxy/G/+un//hvP7x39a+vLoi9HlyRU2YSAHD3B/fvq9kwjhDRbpHcd0Rc6qSmiMg5cxca20/348ef75/eDG/JheRdsEKIxMLtbvcIrUrgInwYy/72ViSVqeScEcndCJEQd7utFRFO6M2qxnLOHHB9sx+GEc0xAB1SSo2abXUF+8MhIhRvrq9vjxLpHyiejNOnTLHrhUWIMQDcwaxLuc9JRByCiCIAkVJKucvqBoiNjg8IZk45A1Lf9V2XmSmcRIRTQocaUTycoCAFsbFMHooILCPRPmAqWszGWvfzrwQsLdDgTh3+S9+Rrys8f0Pu7w053Lf13PuD0MFv60PfsLve/GhfiTfv+e8hB/3uG/9Gn9hGD+6OAES02213u11K3TCML17cHIZR1Ks1C6M7IDqSs+1HOh6w/cXMWkUF3l0rimWwBW3129ogEAgg3Fuya601oIVPBwDNZ7P8j4gJsZSCiAbIDuyBDgiBEI1lJkKECDd3Y3GmQLD2iKNFIg0+hWu4JxYiBIjdduPb2PSSEqfEVxcX3dW9scZzoAmwox/OUuyKFStW/AvCSkCvWLFixTvFB2N6fjVi2j28dxWXu7LrwKZwcwck7Pu+23QQwEg5ZVOvqo3zjeYpEEsJs4WBq5mpAYIildk/gvYL5epmmC8O0Ol0IHAEoKX48UhDu0epehiG1HU555iKmntVc7dw0NoY0Vrr0UYDAAFK+0ub5xCTVlXTFk44q00D3KMR0IDYPKHN7Ghe0U6k1jqOk6rGYp78RThjSOfZzvw6BjQJc9MlN4KYEInDQ01bkjsgEh01O3E8TGOf57gz98U2o22F87YIAOgLwxtLK5aj+Klhd0tTFzvqpiWMcwuPlzDbd5xvgIiITkpISo1hO5HNy2U8iRTjmBQZceLxA9zd1bRWrdVUCRGAIqItRyAiALVTiFmK/V1PzAIAzLxqQaaUs0Ut1ZBgt9t5uEckka5LoNXNhmG4ub6pj0pIun32ghEvLrYXFxdD1NTlzaYjwt3u4jlBKeM4HqRHYSZiiPAy4WHf5J+E9JUt+wK8OYnwNrmSav73Hz/+f//hswc9/buHdJmzBZiZW3g4AGy2W3UbtZR9ee/q4e7yMgCGw2EaD92mf/r0iQUb7W41/+Xf/uPvHr8o+tor+3pJ6hds+U7JIATMOTMmqCU8gMAj2nVUra1KPKeUJTePfFMt0yicc9ddXt4b7z2chnEchntX93e7HdQCplWLDOnp06f97t52d4+QkUjN7l9cPcRtzh9/H/muN8Zo9qKUJ8OY3a/cc+601lqrWSDEyEgY0Qh91TKVUqZmp+3halarCikzq5mZtiWrqnWYRiGekJUwOEXuJhYDOJDs0YrF/jA8PQzPD2NFqO7VbVSt7h6gzQAIAL77J8uKFSsaELHr+pw7CBwO435/cHMFi6jm9tJ3kYgA7hDQS30VAkJ4c7hyJHrlV8BSdAZtnd/asImIIMJCvZYwPcmSX9lZtQxugWQAHCGAEshBjEAICgjgjbymcISQwGAURiJOKSXGTqRPkhMlYSFKSXJq2mcSQWEgDGHocqYuD14o6L3ODiV/F92+YsWKFSu+HCsBvWLFihXvFDvF/+aXD3/672F3eckBlpDRaimlKjF5WLWphfQxsruZWtWqaqZmLc7FvbkqQ4Cautji+BsRDuGhzdjZTBWdnbAT6lo4V1OnHH0kIDxAzYdxTIchgMdhrKpA6BHWlMsAEKFuLeUcCRFo/kSPiGDhlJKqtgr3mIP6MALcwU8EtJtbC1VvFFKEN4a6Vl2S17+y/15HlgXEEkEI8wlio6UDwM3bO0TkQRh+4nAXPt3d28uBGIQvf85CQONxltVef9m44tiGhadrVPhscwHnnhcnEvy05x3q+SgNPFa/Hl8+56AX7rtdpdlSuvHQp2lio/61mqmpOhBiC/w76slhMe54Z0AmEuLQmkQ6QrBSa23RaMKUc2IixDCriJhyAgRwb7cjmCNiQLSTQoSUhRDMVLVyBDEBNoW4R7OCdvNXZF9f2cg/LGPmHs/39ae//OTHDzYfPfjg3pa0lMM4uAMhE+Ht7S0xIwAxd5tNKWUcx1ImxIBw1ULdVfXurz9+/Fe//O3T68OZBPVIJX/RCb5rrvlVzF46iETELAKJCM2diDbb3eW9+8P+VlUPh8MwDgi46Te73QWFA8RwOBxS7xHty9N1mZCKainTOI43Nzfby8ury6s+52msEEGIpqq1Ev9wjFpeB3XfV/18KheEF0laebqZA4R7mDsyttqKVoaiaoEt1zFm3yIA81BTMzFzDzf3YmZmE2FFUEJFMLOitje7VhtDI+LZYbiZihIZuLoXM/XZwdvjzTx+VqxY8TaAiCJ8cbHrur5U3R+GwzA2TYCruttLv+7bc9Ld2oO/KZ0R54KyFiPh4fiaRdyXCWhsFU7EbT8PD5iXw88VBO0XDAGEh4c5zSZpDmGBEBQIhMCIEI7gzRdECBNTSpSENn3e5Nwl6ZNssmw6yUmysAjnnLqcEYMomJAZuA13coJhRIn9eJ/r7Xd9FVasWLFixatYCegVK1aseKf4o6fbX/5xECZ06rouogh7C/dDIgsrOjV2djawUFOtjXxurG6Ee3gTrSHMml/3Rk3PeXqq1hhhzNuCm0c3cbXbMIA2tnZuyzwl0IhxLAg3w1iHYVQzTqm5V7BIALSMGg939+Y0DXGchwSaT1W9OQ1HYCtrb9mD0fhRBECfS+oTERGiuSEAIzcbEFMzrX5uKPEavPJW40zCFhMJiFlwjDEbEIIvtK/N9PTZLGh2NJxFz7gcKM400MctcZZg4xlxfbQxPHJW1KjmY2Njadj5/AtfIvdiPkws+7/iibFM8F7mDQPQlw85tg+ODPri73Emi475jmlq62YFGXfUSe+AKEJETClt+p7CW8hl46kaVd5a4OE6juMweFjuuq7rvRZ3OzqMC3OppZYCCG565O/b9XdXACJhTKmZp399hv28T76SllxWDF7e95sjAKrDr//5yd/99t6f/PGDhxddgJU6ukXOJJynMnlENSXmqqqqwzS56Xa7ifDc9cqb3z8Z/tNf/u0//vPTw1Tj5cN/r9Hs49vTDTGYKTyqFndHgtzl5kpUSim1QvOpEW6G8hGhVo9W4M08Z6ZZIWqt93Pf9z0SlVoDgJgCwt2WFaM3bSMA/MGZ+pdQIj6t+sGmSyl1XTd6RACxpJRz6jDcwCUlYo6lpMPMEFGSdH1PzA6g5i0z0AMDKYiVqCCOEWNVNcdap1pvx+F2bPZMcjuVQRVSsubwHmHu7fH7vb/XVqz4FwVmyjk/ePBgs93sh/3tYT+ViTg54Bf9Jgx3aEZpgLFYqc0r34wRgT7z1Hf2OlpwLEvsBMCNLUagwBoW4TAHGM6jlbOVdmTixNwlyYHJHc3QHWefkBBERkxEOacuSc4sjDlRl6nvuk2Xt13KjIkxCTI7oxMq1jLW2ySUk0ifO0mSuHp4ZmCIIHj82P7oj77DC7BixYoVK74AKwG9YsWKFe8U+Gd/9hf/x//s4/Dp577bbKlcC1ZmIhZOAggWs76RmQ0wPEQSS0LEVsd8riJpMeJNiezuR3+ICHC3UmpwN0X34fv+8N5Fh2AAfqJWG9MZGGBm/Wbz4Y9+fHNzexhGD7cAQJCcmlAOmQJC1eYZSJz0ts3bIhaqgZmJ5lg/d/C52BOPetJmajwTgh6AkHNm5v3tzTgMPovlvpyxOPGwL+UFYkAsIX5xtuVMtiLE2fTprt/Ekip4/OOcgAacwwnbwWPhfJuvxumYZ4XmJ27qTvYhwilz8NSOuTHhgHdfPmvCy3+NOUj+rlr7dT4mcfxn9i45pg7OLTt5Un+VMPbtABFEWHLilHyMqY7kNbEQUilq7uqGonW/L8NQSqHw3HduXkvBnIlZmHNKVrVdqmkaAYNwDseMcHcNTCAEzJLS0dTyazXz62/8lvstAJ7ejL/4zec/+1f3Pnr4xw84ScpBLpK6bgMUh/1NqTV13c3N7Wa7bQ8KFtHwzfbB71/AX/3yd//pL//m+b7Yy4L7lz7nta+/hHfNtP5/7L1JjyRJlib2NhFVW9zDIzJyqezaeqq7ulk9vQ67Z0hwgJnrHHmYn8EbeSNQV55544UgQIAgeOOVINgggQHB7qrh9MZau7OqOveMxRczUxV5Cw+iZu4ee2ZGZkRG6YfMcHN1XcVURUW+973vtV7FvEY4EXqYaq1ahu3FuF0RkbAAMxEHQq11t92WUpfLbrVadV3a7OMOrfZgSqnr+r5fdF2n6lW9mlfT1gmyMKf86ETxx+Llop4biseHpX5bDSDU1NSgkestg8a0lKpVI4KI2kPfyglU9e04MouwFOedgzoAACAASURBVI8EWBFNWEOC2AM3Zqdj2XoooCM0r+fBvQICQAVUQK/VWiJD+CE49mX6y8+Y8euMZkEmIsvl8ubNm13uTk/PSikAKEkCyK9F4a9t6sYxpYtxGxS08oQRERyPzgjap3jBNJpqumkChAh3M2i89kPb4t7DjBGFmALRHT0EsY0NiCARZqIslIS7lJJwK0ucBfucmFEoMMw9agQERiAyEktLsmMmSSLMgOiB0veFpQB5OPyrfwXvvPPcG3/GjBkzZjwVMwE9Y8aMGV82ai0Q+MlwVmslPWMbE1NKSVJCJodgJhHpUjIzN4/wVnbQceKXCRGJGvFJMI36W1Y1RHh4KzOlWg1SjvTmbb59crRgGOxaKvRBzFK1ppy//vWv37t3//zioqpWMw8nYfdQVRIGANWmM51ozIjAiL0+eJqFEFEjaz3APSbzzzalAXAzIiJmgLB96b8kIiymtdYSxZ6JrdgnjB9+v6Rx9xzsoWYjTCJgB3zQgfmyNa7xhw+6cDTmeH+tGOGtyDtcsf64vl+4JPUuzzMumZjLH3s1NbSJ3qOWw/WzjAONHdeZ8sPGB4HR4dPhwHhFGv0Aqx0Hc5Yv2n0iIoZx3Gx3kVI1zRHCzMymvrnYBCIxg0OStF6v73wEZ2enu91u/eYJpwQArrrbbOtuXC2WR0dHgGCmGODhANF1aUOeUkKAYbMx+9iVPr38+WXhFtXhnQ/v/+AnH/zT7377+DV5/fW1jnWzGZnE0ZkEotRS+sUySVeKlzrGWNY3TiIfv/PR+z/40T9+eDo+20P10gERVTUoRGSx7MKSo56dlbHsLjbn2+3O3ftFz0y1FEIaxxKqiTkLt4fe3cdhcLjPhJzTDqCUAiFMebFcH53cUKvmuhutG8dxjLHUL9eL5vmjRNypem6uEVW1udvvsyDA1GtVnWquCgIhBiEFmJpvS5EUCVERBHAAHJEGJAhQszO101K2FhXQwqt7da8BhoAeFUAhVLX5GUVcCSTig3ZFADDromc8J8w30gFTU6SUlsvl0dERMd2/f1+rMnPOOQAdkB9yckbYF2qOAEQmjABz5z0BzUzuzXnt8lhTGYq9LjoACJwJpxiwWYSF+yMziBCAAAkxkXQkCUMAGSMRZeEuSWJKzIkoJ8rCKTX2GSg0MXU5Axq2wofmji27hYkEpyFQBJIHlmqghswpLTalbAwKKL3zH/jbf/jFfhUzZsyYMeNRmAnoGTNmzPiyoRHo1SAwIYOA7nQsNu6IOQDcXd2IadEviWjvZRHN+tnMqio3gTSSMAsLEaWUck6t0F+TIhORiAgnof5NWb158+jGEjY72NXGmjZ7VYwIi9juht1uW7WYV8RYLHKH4BFVzdyJsQlIRahNJ1ikTSh4ym2PlDIhx96guk1m3GJP+aIkacUM2+VUrYiQEqtqQBADC4uI1ToZOl/jVR+ZMoqTAhwOhO+h3l9T+zZO+iASbrLtx8g/H7H8yl+h2Uw3lc1+eTx527jy82FnhgeuaGLJn4b9TO5aEz2wT7x66Ad2+cCCRzbrU0/i0+PBL9QdzEJNrVZi7vOCdNwMY079rVu37ty9s90Nb7x1LKnb3L3r5uv1Ud91WDUxQ4Sp5q4rFz6FZwA4pdT3HWFOebfb1qpmxk7M3C2X+vE5THWWnh1XRcGPmkA/6Uqv7uHzIgDOt/Uf3jv7yx9/8Poffa2PIlYJYdgNqZPVatUtuqoKEZuLCxK5cXKSFpn7G3eG9JP37v/0lx8+g6r3ZWHbryIimvE9Mo9ld+/uvSRyenZvu9um1OXUE21VbdiNpVREIpbjoxu7s9Pdbnv33p3lammqIrxcLvr10TiO43a73W0DYLVcQfg47rab891ugwQiEgAWzswv+ro/LzxiZ34RsQFc7R3kU065yymlMEVCYmKRlEREtJneIAYRSnJOlcWQR6Jz9zPzbVVTK6QX5hfVdu4V0AGqe1Ur7hqBhNVNDwkscegcG+Kx3fiMGZ8R8x31WHRdd7ReC1EZxvun9z28y7nLGYgBEenBHn+K08P0rsM2EFWj5piGhDQVuYZDKeaIiKhm+1wKAIgwJyIhKnUspRUkoQAHf/CbIsSMlFnWXX+UsoRnAEEQCCYUQiYgQmSw8KJuYSIkjIJBEdWNmVgYmZiQWs0RJmOxiNAwi20ZIYY67gCBcyebUkgKioLAxf3/5vvf/+K/hxkzZsyY8SBmAnrGjBkzvnSQKWcftmOtLdHR3UK1KVo9wiGQGGIq1rfX8EatpVZVVRFhYULKKSVJTSdopm4eENjmCohEFOgG5tAntGUHaQQC8OsGFhFRSr242Ny/f+/s7Gw3DCwy8QhIPpl7NFFzM3o+uCdDThkAzKxwaXaB3uyoWxa2BdFU1IuYAcBUASAAqmpAIGIptVWrUtXLAoHPpMDdl1KctNeHKRRc3/YhDvZxe7uGhx0VHsn2Pnyqj05u/ZRHfwIe55bw1EM8mWH/0t0VJuNzkCRMZiXGcSTiJAkAEKjvFwBgZsTUSyIirdXMIKKqmqqpGTeHgQiIcRwDIaWUiJkJCRGRRGS5JNlOTtOf8WQ/W+M8NxW5Wnx8/+Iv/+4ffv9bN2+kdENQIKzWqC6pR+SiY9f37oHoOUu/PNp49//94qO/+em7739y9mlrL75MCCYmYXLGIPdAkr5bLldHi8Vq2w+SOiRGoPZVM3EjTIgwp1RyAiKLMAck7vo8juLnNg67G4ueQt0GREeE1l0iOrycZPynQQBYxGnRD4bx1tFRM0B3s/Bo6fGA6BFqVlQ13AAcUQEVUZEcMQJGVfYQ8/vDuCvFEUfinfnGfHSvAY6g5tW0ejgEOFjz7J4CfY88rwfxhF5sxowZnxYHB671ev3GG2+KpIuL07t377obM9dagRyI8FEvwweyw1oJEroEItI17rmpjz0cApvF897jS92mF7T7XiZ9+bTH/lSBMDXffiK2QAjch6/M91sBEoIhMLgBWaBhuKOFMxMbKzNhAHi4iXDO+VBikQAIIsyAiA3KqIXBEyniw4T4jBkzZsz4cjAT0DNmzJjxZSMQOhq3AVYUF8LMbmSIbuYRgUDCxOzhqhbhCMjMSDSWUksxd0CYaOBJqxKllHFkN2vl3cwtIkTEHKtTpYXV3aqntGmj/AfPqGrdbLd37tw5Pz8fhiEIGxfcLReAqBYR7ubmNrHMU1FEWCwWhFQn7hiJqOmfoc1MHGhf1Csmp+pgJiTyfUWwWmv7WMdi9mBx9mdozQCYSPrDts+DQnrCaVyleh9JMn5+lvmpOMzn8KHlj8SzN8kXZ75xbc9TiTkkQDQzVQ33WouaCafcASAAE7M0x3DzvXmLO0xxDosIJAQiIqxa3b3r+9QvRAQAzN3cGyuNiC9ixvl8GjMANkP5yTsf/uiXd95av74+SRmK14qAOpRqFuaMCGjRkiAwfXKhf/E3f/93f//uxbZ8/hN4IWhBJWJumQvEIkSJu8RdlxfMSTgnySjCLABASO2WkJSXy2XOGQCqaimFcwWElHNKEhGqVYTCq9YxvHoo80KEifyr7r9xwL1S/nGz+63bIIjm3mrS+t4Wo5qPte7KOJoFYgUsAGPALsA8NOxiNzgAMZ/vhqIaRJVscNi6V3ONcAB1q2a+74J9X93sGVvwwXJmDa/MFzBjxgtBBAIcr4++9tZbwrLdbu/euavmgLAbBkAC4n2xiqsbPfjYRUSEIx7oZ8Crz/iBhW7srxkc3tgICKCqqtWsgj8iIBUABuEQjQwPCPVWecQJ0RGIwCCY0ByZkBgNkMPVgNErgSgRIREJE7iFKYSnlPq+d6+IIJIYIRH1KWESSB3kpAEWbuG5fmHtP2PGjBkznoiZgJ4xY8aMLxum6oJdSjdO1m/ePIHdArS4WdVazdQDm2g4XKuqajNKDoTUd5RShCdJRNSEyVVdaz3MCloWJRIBgJkFclBSGCn8zdu339uc8XbQRhgANK+KAFB1VQ8Hkdz1+6p6iJJTBCKaRxg5mDWxIIg0PplIkDAhNa3LnoYAYmZsWd3UlDU2UWPeigRaTBXvRCTCVQ0gPB4p1nwUI/Eg7xpXWeEnbf8I0d0zcbiPWenJbMkXyqV8zp0fuNEvU/F5eaypbCaiVh3qgG65y2en5xHR9V1UrLVg33FOETHWWktdnfSLaqGVCZNIRDCzpISJc04pCbszc9Pgq1pE6DDqZjMlCE8uKl8yHnZf+SyoFvfOxx/86FffeG352vrWLWFw5462m42a96tFGXYGZoBV+mHnP/7V/R/+3Tu/+uDOV1f+vHdtQFWPUompX63CwtxrsTJUVXP3hEBEkxdOgLkDYM5ZVbfb7bDbqWqEaymBYepMslgszHwoFcZSSlW1JCIiSPpIUvRppwkvoWz6XO2DsQ4Wq8AWuSEmRHDw6m6AFbkAF6DqgFU3Vc/GelZqQa2Am1I9AhA3Y6nuwGwYJWJQre7m4BAW7h4OfvkuORz+of758i/7Jj6UDoiDNVAANL/qw3azJnrGg7h81T+fvvUVAyIE5Jz6vh/G4fT09O69u5wykiSWJhVWN79OCk+lO67tBlu1EZjoZtgXGbnOQTddgXk7MgISI13b1ZV+4UpeGSIiYRCOoVENxpIwMiEBMgI7ICIbMCERkiITIgSCM4cwCAMhMmJiZATGEKREmAgAKQn1fWYMIVx0KYhdxLtUq6HDySkM/RfU+jNmzJgx4ymYCegZM2bM+LKhFrrz28fLLqW+6916SoIIZlbda8tjjkB0V2vi0KYRPoCZIaLW6uquTkThcVABm3szIGgCQmARTLdOjr79za//7ON38O6AiHDVPHnPBpo5BCDQNDmJ0Goe0ExCPcIjCLBpr9tURM3JJ7aaAAMAgQJ9SsOetC97cmHybMbDckIiQjMAMMBHS+KunObTgFcO9ax4MnN0kFQ/uNoji2o9ctuXGC+CjwWAPdFELCEJACIgSbpxfKMOGuHDsC2mCADbHVQl4iDbDWU5jmf37xHi8XpVxgJAYynb83NMWbV2KTMGEdVazs5OAWGxXC4XS/cYNlur+iwe2y8zqvt/+PEv/snbt79262h9W27cuHF2fkHMfUpuPoxjt+jON9thi15u/u//7q9//suPt0P9al9zACKulisRgBo6FiHabrbbi+3JcRDibrcrWk1LSoKIkgQgdrvt2dlp1/XDMJoZIwngarEsu40gd3lxevrertLq9a8dn7yxXNVf/sOvLs7PF+ubXc7M/Iiaol9BbM3vlnpvGAEpABzQADS8mI1uSjw6XKhtHQazYTduq16Ucq4+QpSAbVGHCMTBXc2bGFIdipl684naM1BTQdQndiXtFdGq1DYr2en9NGXwxBWnqWg+s4ifSk8941XEk8YD+LyCe68WiKjPXd8vWGTYDZvNdhhKciAOQG7+PJMzxlVEPDohYf+hma414hkmrUNERNDVoDK4mwECoh8O0R7ya8WvL3dibqW6e2CtwETIHE25ANRMOCLaEnBECMJo0cZAQERmZKLMlIU64S6lvktMmBP3fSIMoehEIGXIy00QeAmDYVn7bXqejT5jxowZM54ZMwE9Y8aMGV82tMTNVccIdRzLOHoZGSKlJKljggSgpgCRk9DkEO1NB91qBro7AJjZuBvqWBU1WJhIRKaigu64L0KIxECM0jl3ZyP8xU8/Ibw3zf3jmoWEe7SjqNaiui9mSA5h0MxDMSIYudEHZubuQtZ475y7lsFOiAikqm7hPlWnmawSAMId9vVqEFu19DbL8HbCpg8ThQ/bMT8ez4FTfTb76Qc/PC98mov9qh4R9pESm7gowvAotZqbm6eUpetSTiBCzBiAJMdHRyTSmH8ESCKI2OXcLxbSZXUd60ju/WJ1dPOmue4uTs0diKjrht0dM/9MxGI8LUTx5G3h02/+2NsvAs629tc/e/9brx998+Tt3sfULYbdoGb9arlM67und4PzEN2PfvbeX/7Nz++ebb7SRpeIKJIoZ4udRAhjqBPRcrlar4/6xUKtLpeLwDC33bDbbDe1VGZBhGEY1uvjGzdOdKzb7dbdN+fnBN5Uk0fro7xa5dwDECCmlAixqm42utsNz2wCgZ/v9vhiUdzPan3/4iJE1D3CyX2nujMdPSrx1t12w6nqtirEZvAY1LcOJWL02GqrNksFSCFczQHco7p7gF+RNT5zY02kMxHSXlrZ/jNs+sqpPb1x0IiN435hUbIZLxj40j5cLzOE5eTkZLVaAeJ2txuGAYFqtagRgIAYiA+7sPmjjDIA4CAiAID2EB82mNLnRJAZ9zlGZhFmBlM1agAAIsAAi2ujJowIMPMaFcI9XACCBOCyBuzBuw2juTkjETJjJ5AypkSZJYskokWWRZY+SRZJwn2fc2KiYHKiYADpl7Q63p5tWieDgd//8z9/Ho09Y8aMGTM+NWYCesaMGTO+bPyb/+K//Yv//r9k2JWtnvGdzd2PwCszIyEygTARCXMSCfdwB4DJhm8akAcLE2JOSZA9BSIQETMjEkCYe3gb7mPTUoNZJ3L71s1ln4Um/uBgItw8+CJctd68eZJyOrvYNDtmB7RwNSNiJEJAJkYi2Fe1SiwA4O7M7RQIADxCVd28EYBtBSIMAHNHRER0N0QkZkRw86JVq4674fT+/XEcVPW6vOlh2+rP2vrPuuGjskav4zMQtwjSfAI+zUZP3N8jljxmGvngVg9w6F82yRMB4QFqZsYR4V5LMZ2qHgUCi2DOjYoSkpQzRiwWfbN2bhorJm7+zqUUN6vjOI7DjclygE11GMc+QpIQ0zOc1PPlOx5o52dh0p6yTnX4h/fv/M3ff/Ddt24sX+fVsiczc6MkhpgX6+L5k4/LX/7tL9796HQo+vmv4cWi5XSbmVllZMAw07Y8wmotSMGMzBjR0j5aX8Rd1wFA67UCgJjUjNGr1qEOzJiECMx01FqYcBxLKmVvkvyMeNl50Rrx0Vg64uOuUxYirpIG4h3iiFjdN6Wcqu3MAGk0H1S3pZaIGj6aGYCbmqm1NPtJ4eh+Jc9k31qPsy2aHihCEOGWFMMICIERjMhESNwqi7JIS8PRAAeY2GeEKWPmS2iv54Bn6UC+/Et5jt3as8dmnrqHxoJetVs5RHT2RGdECxG1z5c7verkAM/97vj81/ip1nn2Iz79MIiYhNer1froqO/7+6f3N9vNer1GEiAKQGvFPRABr/k+T3Ya3rTRAQDMLMLtb4fVPK4poKF9i4g4DTUjIpiQsXlAq6lHo6qv9BnteWaAjLiS1CF0CAkwMydmAmAAwiBAhhCEJJSYhUkYmbHLkBOIYM65S6lPOTMnpi4lISREYY6IUhUpCJ0whBVLPRvGQX151ql8dY2pZsyYMeMrj5mAnjFjxowXgPBy4d2aah2wjLs6DtGUJowozEzMnIjd3M2JMKWUcwbAgHB3SYmZEagN/wkJEGOfJsnMPlWL2U/Nwhc53b518+R4tejTZquHORvu/zHT3bD95vFv3Dg54bv3TJvtBqi7qiJRBJi6yFQUbk9AMwBY84aeSHCMCGVuMxkmBgR3b1MUc0OiJqAGAGIiRPdgE0tGiLvtptYKoI/i714InixyxGfw4ri68sH75DPj0CyfR5n7TLbXXxz2tFVErUk4UYLwQJQkHmGmQRjhQKim4Y5JICDUGCm40RMRHoiIEKZqZiKi41iGoey2WisRIaG7gdliuWDhl0BO92R++ennFwD3zrc//uVHf/XWybdvf2fBiVKy6mNVlJyWJ2WDv/z49K9+8qvtYF9p+TMAQIC7gzsxAkaA5ZS2YeNYdsO21NFcax0ydcwsIqnLyFxrRYT1+ngYxt12O4yjmQNRWvRRRzWrtdQ6iGZwBVerxU3HYexUifacyysB9fhwGBcsi8VSAap7mJ+Zn5sXh6gaEferjmYeUM2L6rbWGq4B6m4RFh4+lcaFFjSKy9vqyRLolrLfntUWWsVADCAECkCIzCwsxNwqnS1XSzcbx7IpQ/OfBghwcMCviAr62RW7rzwH/XRjq8mKa/9rACLEVCk2sC3dj1L2g5Trb9qJ9dz/7VNcwdPxLJHC5/s6eT4cNAIw83q9Xi2XInJ6dnax2aScWDKSOECjhJFbLxcHDtqj1a8lc3cPABDmnK/5VEyPf+y3jGuh6+bJAQCNgA4PB/WJlr5K+AYEEIAAdEQLlgVTh5gBmIgJGYAAEIIBhDAz5sQ5SRJOjCLYd5gEmCKllFNepNxiFEyEAOE+jmahVStxEAWEixM6X+zGgpIA5OYnn7O1Z8yYMWPGZ8ZMQM+YMWPGC8DJJp119/P6aLla9PLG9vz+sNsBhIZX1WGobs6I4AEBTCQppSREbGZDGZmZqA3XiYCYGAgBsQk/mxfHVLycGJGYeLXo3+y7r71x+7WT43vDPbNoRpuHUyql3Lt7N6V08+bNsaiZAaE5mE0eoMMw7rZn5p5EEEnVrKqJNDU0cit76M3xz/b0V6OkAcDdW1omEiFANQ0AImqqm8ZHl1os4uH80BeBq3Pax7K98eCaT0b407XPnyr9/1MhHvr8VJ3aF/FN7AMlbcZrenLjhHU7XoDVckSy2WzGUnKfaxl93NVxV+pA1AGCm52fnUmSkxs3EJGYkNDNQ7Xv+rHv0RQJt9utmkVE1/Wr1QqRhOWQQPAQ8IFze97Xi0/8Fa409QNt/ujvtxr88qPTH/70/X/xR99LRQWhWt2V+sZvvHZvh+/e2/7svbNffXC3+isg8orwAPdu2Qn0ZNb3/cXFZqzjMGwjbL1eqioxA0BTOpt71SoswulsONvstsMwaHXTWK7WZRtJODHVMmYtQpiFR/CxVBEWYaw41at8JaDuH2x3HeIxcwmISqJlMwybcSwWUdWZz8dS3AzRHNRsrGrNJTaiWT3HvgIZwKVk8lmiKO1FMNUlAwhzYUyECEAOhLDIOUlmJGBfLPq333qzqp6enb9/5+PtWAMJAypGBcCIZzHdn/GVwlVPBkAIBJD2ZgAHAAdQiEku35ZPjDPuP803xIPwCGQ+Oj7OXVdKubjYnF9sazEJIoEAKLWau6RAxKmAYIAfyOM9IkLNolzbOcIVB46Y7HEOlTsQoRUXCfdqVms1VXe7on2+titBzIiZMAEkAI6gCIpJ/d72SUS5y13iLJITi1ASWPYsDOFGgGFRQcPNzbFpH8KGcaxWgSInZgbVktdGCmN1J4R/9efwzre/oPafMWPGjBlPxUxAz5gxY8YLwKrEb999+29/ZxtI6+Nbi76vpgDhbmp1HMdai6uampsdajFFgEWouQcQBqE3azxDRpwKuzUPzUZACzNSKxXOIYsqqz7z0WqR8H6Ax3WOVc22w/j++x+Zw/n5RalVzQGpWX+qNU+OKHXcwTglYHrE/vMkfFYFRELEy9I004dDwSoiAoSx1ojAfbEadwNAN7PPTjN8GurwSfxtPOzu+tDs6eH1n2XP7e/YZNNPu86rk/OrRzxor/wLS0x/OvP+ufcMHs2PBYZxt6QQJnfb7TaTQaUFmNezM2rcIiKnFBYeNo467BIRIGJzLRciANhtdzYWkYTM3sSbEUQMfVfreYQ/gwX0Cwl9PPCkHNr80XdSAJxu69/96u7/9u9//p9+d/2d1+Xm8ZHwArH/4P7F//nDH/9ff/HjzU5fBbZuijHQJMkD2mx3iHjz5OTmrddXy9Undz5eL9fWaqVanJ6e73YDS+eA733w/rd/67f6Re9qZ6fnfdd5KeguTIlFiI5XawzcnG8vzjemenx8IizDZrPZbOMrLx2f4BGbWu+N5aM0AhEyE8LOfOs+mnlEmG1Uq7sDekxVcD3CWngIWq3Ba14b8Kib8oHuqXVYe3d3JGgWrpCQMhMDMEVCPFks18vVsu8Jabno33z99YvNhqpuUiYHQwJAB2uSS58LEr4imExV8Ep/15YK4brDb7z99je+/hu/+NW7H3xy997Z1ts4A1pYaDIvbh4OAXsJ9HxbXGmDLOnWrVs55812t9ntSikA7O5htpcjT/H+Q1HrNgKLgGnY1lJPENwc4PLxRrisUxgx6dMfjK8GQHi4mao38w18MEyPewJaEBmBmrNPK29CSERMJESBGMxOXIHco1Znc1EYVQk9TCGCEIQoXN01wpkwMTs4IgoRECGicBZK7sEQ5rH90XeXv/uTL+x7mDFjxowZT8FMQM+YMWPGC8DbF0c///pgQdviN9bLrs/AjZV0cK211lLKuNOqplprbRX/ABAqqTe3U8QA9EAPBJ8MFCPMfBwLABIhESERIHpgpF5zyYLHqy4h1n1+6yGLMjyq63vvfbDZ7AJhtxvGsSAzIAFiqUosq9VKVatW9xBiJlatzQkBENrEJgCIsKmwoUmho7kONkyu0GMpthdpTlMPwDYN+kzTyU+TEotX/o2HlsNE5j9t+6s/9+s/Rb2Kh/+bpO8qr/PQpofsYry664M+PNpuLnfwaZvtRZGtU8K1mY3juNlubxyhuw3jOA6jux8fHyNeRETf9wDgZojIIpAzAnXLpZXRXUutpRazBRBT7nwYGuGVJK3XRxFRtuduXoaBtjsKukzX/lz4IiTST8WDTLR5fHx68X/8P3/9xvE/vX1066gTCBoL/vufvPtXP3nvgzvn9qowMggYEYjk5jZWIgSAYdhtthfH9YaqIlJmQsAyjMJytDqKnBGROZ3du7/dbNyMCRFi2G4pFCKIqO96LeYaWfJ6sc7S7bZbWRzlLl8+Xc+ELy5R4Dkg9qUIPxyGnFNCIKPBfecxmLmHE+3UzB2Q2rujvWb8SnL+U2X5DwbHpuqC0SKfREQRBEAIHXMvkgg7xJ75jeOjm0fHR+sjDMg53Votk9Yt83FK6FGJ1UO9MV1NEjtz0K8Grr16D2/jTujNm6t/9nvf+bP/+J/933/xw7/6u5/uNrvioeE4WVfhwYkDr1pyfDUcWr5AHK5eiBd9/9prr0nKd+/d3e2GqirC5g4BgdCCeao2Df8mQEo45QAAIABJREFUJ40w87hSMro9/Y7TCA0fH7y9Nl5ro5MIiKaceGwWDgJwI6ABMDya9TREIJIwg0Qz7fHAamjeeHFGYAIGh9AwhXDCEEIEB9AITUkWXdd1ucuSk+QsiZkCUrcawoRYXe1s9f3vf67WnjFjxowZnwczAT1jxowZLwD4/e//8H/8r8LidLNbpAuwneuIGMxEzMxMCCnlnPKVki9Q1VppF2bGVpCrqqkSQPhBz+KLhU2Kln1+pZo5BKEfrxcn6xUTXiUUJooBgRDc1VxT7kS4FGjuzyyJiCJ8s9moqrkTcggEg7cs7eb4F9B00KYRbsRESG4BEMSEiESTMwgAEFNL+2Rm2Atz3K6qfZ8yp2zHevYmh32i6AM7ufrL4Sce/rAnjSft8gPbtM8T6XJ913vdz3XCG/YMLEyu349A+KUNSWNzcNokIny6IzwswqYm2E8jHzz8k/C4FR7pEfEcKbYpVICIhITNORxsKmGZMzF7TJNh6XsSaTfNJBv3iAgiWiyWOeWu71PfAXPVight6hlxsHuJ8EAzM28T7Me3wzNe4BdKNT7uG3lweQDsiv783U/+9p07XztZdpISjh+Pp3/1s/d++dH9XX0FzDcaJhOH1vshobBUKONYttvtOI4ppVorEYWHSFr2/f37Omw3qeuOb73GSKEG7uAxDjs3i1AzQ4T1eqXmbiYsy8WSEB1ARFIiEXlpCeXPhq3ZB+Nwg6gnRqhD1aHqoObggNQkz1PCgEeL/01y4yshmyfxzvv+ECMQkScCGgVBmLJImEGEEK5TPl4s1l1ed+k459s3Tlb9goE/+eTjs3FIu43V2ntdE0KWylJqVZ1S8cO9ndWvPdn4SuFwFwnAjeXyn//x7//pH/7ud7/1Jup/RFE//vD908F3Cq1CQAAeTMOivUNmLw4AgGjPXEQslouTmzdvv/baUMZ79+4Nw6BmyO7F3MER2khMzaLZmyDsZQEY+54W9nKBRx4Mr/TJ8NAICgMAzD0gHMIf99VMg4CIpswOcwiLFmZwB9DJBhqBiREDEYQoCSchDKMwDCdGYQThvktd1wujMInwou/6LvVJhIgZExAtFsN2gwBTTt+MGTNmzHhxmAnoGTNmzHgxaGyYAziDVdttz8MKQCCziAgJATIhAQYEIiJSeGCENI6aCISTiKu526VuduIiEWDvbtGIOM4qq7ffeO2N1+4lIoLrbsRT0jSoVrea0hIgA0apCsgkIj4dIQl7ACGJCDPHntdz9zalaSTGNK8hFGEEQAJonKMwEkEEIphPPOMkoDYzMxHGCG/ugY/llxshi4iTPvjALu95bpwOj3iNI4Y9O4KISMwEgBGO+121VabpLRw23Iu3WwvvC3G1fNXDOleI4mkxTJO0KxLmy8VTtGC6nsuTm7SHE4EKgQfJc4RHuE1fqbm6qzdu1fx6kvrnnJA/QPJ8IXwcM/d9t+gXiDUAhKXv+3EYaqm1VCSMCM5dypkITRVqDYsyDACeUko5LxfL3Peckk/fFna5SyLb7Xa73ZRSupxSzpiz6sVBif+Y630Z8DC39li2zQN2Jf7qpx/cPl4BSMfx0w8//MmvPrp/Mbw6ZEyEu18+hUTEZDbFKgCCmbXW9rDklAfajcP27PRev1y//jVZH623p/cR0N20FGYKRwSk/eMYV+R7OWdmRgzmT1WE8CW5c56E6n5RFbgMEUxUVEvValN2fXOq2Qex9p1P2/KhOwmvL2oXT1MwCSGCABK3YBEIQGZZ5C7MEvNqsThZr24s+gVjh7BAPEmpZwoHrmMZtjR2ya13PRJmpkKyE65mGAjmAeABDjHbQb9KOKia/8k3v/Ynv/edf/0v//Q3v/7W8Wrxe9/91qLj9bL7wd/8/Ge//PDetujUFdCeg97LqH+NbwVC2j+y0CLUi8Xi+Mbxar06/3Bz587dUioAtEoJFs2bDYH2YoXGXNM0KjqYOMM+un+QQl9BTOOZ5n2y7y0u4/UtuwuvlId83MmTIIl5gDuGR3MUw2lkjBDUhngMREAEhCgUiTGzMDKBi1BKkpN0mXOWLCxMTCTCWTiLYHORzh3lnseRq0qhUX+N75gZM2bMeAkwE9AzZsyY8WKAiI6EiJI5ItdzHYeN6mjhjMzICRJPLhZGRCLSOF8ATClJEm5FBhPX6gBA+3J/AJBSZmLflywXluBcsf9G4a/96l7mByttHXwhqha1kjvJneQulaoOAMiNZCBqwhSEAGImpHDfT0X2kut21L0ml5jarKLZDnKSNrfpcvKIZjLYSOMmW8UAjCjjGPFEN449pX31qomIiVkaP08siZgbDY0AuOelA4CYRCSljIhmRk0JNDHX0DTdcFDp0kR/7WljV9WIdmmX3+aB5A5spZP2wYC45McPFLM36fghh3hizukwn27uxu4OLdM4JpmimzeYq2nRWmqpCmoaV+Tsnx/PUWj4iDkoAghTziklMRvGiwsfdgiwudisj9YsPJGMpRCAmYUZlOKBEI197i7u3a1a6zDoMKa+P1otd4kDwtwNYBwHrUrEedHXfhFXCxs9/qxeAjx8Vo89Twf48S8+XvSLbcWjXv7fH//iF+/f3476hZ7flwl3L6U4QNf3US52m41LGoehX/Q3T06Wy+Unn3zSiq4S4zBuz89Ou5xvHB8H4Om9u8uuP3itHx0diTBjTwDjWP7x3ffefPNtIqpax1Jy141lrKW2nmuf6P+ir/85wSOK2fkw7KomZvNQt/Cpj5vstfdU/GW8DKbFh4/Xab/JbYNar9scV8MJomNmJApkjEVO625BEIu+f+O1268dr4+6BOPg240Pg5QiiIGUwgNjLTRWreE3kmSggXiTUjWnQASLACOACAeI8JmD/krjamCWEBPRn/7hd//zf/Mv/+QPvsdhp/fufvvrb3z7m2//iz/74//hf/pfN9t/t333bhtfGMIVDrrhcEv+emEaMITblcBzv+iPjo8l590w3Ll7t5oSkzC2gRUEISEQEtAh8NR21XxNWKZ0NCJyc1U99AzT0KWVDtlX+Ig4CNMPYyEkwgBqf5iMUiZKOq6ePUtCElXzCPSIAIymdQZCQAJGSkxdSsKQGHPmPnGfZbVIWZDAWmnuLknTIXRZEjEhmStCUFNgEFLKmBKABPq9e9H3L+erf8aMGTN+XTAT0DNmzJjxYrChzUmsg5MD9svlyc0TWyazGhiMTMHoaKXWsSppeLj5qGOb+0cEIrDIQbiLSM15GQDNjAgRCRAbiZkloXRGC1fNBD2CIJSAuDKPb1qWYTcOiyLCzCwsXY/qbu7RiGLi2DPGbSsigQiPIGTBvcAYwM2h5XV6AAISjMOopojILETk4ea2FxEjNQbazM2QSJK4q/njGdUI2JO5cGCKkdrUqF3LXr/jTSuNDogRiO6GRs1TW0Ta5CsgwCdROAIQEk/Udrj73u5jzyQTIVzlNPHgz3H1jKeU0ksaJ/AgM7wuLQoIAmiCdYCW4no4l+lAbRHuJ4BEwjTNHN2b60RAXJ1cfX4d9OfEI/eAVz+5u2QZVMdhl5kQse97rRoQLOxa3LXr+0Siqpz7plR1s4uLi+12s1qtOIlF3L9/f7fdLXJi5pT7ruts0VXVs/v3cyyEpnn187u0lwIW8NN//OhsNx6vFj9754Pzob5KNAwSCif0KKWC1hZ46/vF3bv3iGS5PtrthgjXWss4Wq3b3YUAdv0CADKFjRuvBcKJqAXktpuzzcVZGcfbr91iYWHuchcB4zgerddd19n5NjxekZvjOsw9QCdz50luuCeuDt3T9ONqBwZw5Wk5pIEgALUCYoiZKBEzUbghRC8sgAlpvVjcOjq6fXITwgWp77reDbalbM59N6Bq5NxYtOROxOucOgJUhSiZ01G/HFUdQNQR0QG8emnuQ7+GdOOrBWzx7gAGeOvW0R9/71v//A9+6+uv37y4+zGYWh1OxwsSIVl8662b3/vNr9/5+PxetQpACAZgPllwTA4cv5a3Q1xa5uBBiXx8fHx8fHxxcbHb7Zh5tVpVVRFJHQAgICMRAPgUAfcW+yZC92uGYPsBSneZ+NVceRCn+HcbFAbkTkQus0YwwFW1lsHVdZ/Edj1egIAIBA4RbqoRxgAswsg8GccDIwhBZswimTEJdZk7oS5RYkiCSVJKWYSFMImkJF3OTAQBpQweDoRmUzHEOgxb16J+cgL377+SHfyMGTNmfGUwE9AzZsyY8WKgWH4kP/9e+j1379brhMde2F0DkJEwEAx0rJqruamqqXm4qVVVM/UI3muOG1UaAK303969ARBRa1VVISbpIY2geZnp1nF3VsputEtPzcltFdVsHEspJaUuHCzczNRskgVOklxkkla1nIgbRTu5WjS1cUAjbSnIzBGDGKupqhKRmSORTlJeg0kZTDFNaxoxDdM5PWlqeS0bu9laNKdQ8jAk8kBSbET43uQiANwMEJhZzUVkP4edjDEAgQAb/47UiivGVZ+PdjCAmNjzvfa5rTNltgLuZcuX6zdnkogm49tTP/t9XiqMYJqd74vIH9jtyYQjwNtUEImIhMhatUl0j2un+BLKOC/nfkTIjOFey0jCqctotlgstNZh2HESIi6llGGwUlPHSGSm7o4QWisRm4aqeVWotbWVqZpq6jmlJJJawIFJRKSFTF625viccIDz7VjtXk4XZ7vyaI/rryyYuOs6rbrb7aQaEwWAmhJRRJRScs4iyd0inNBv3bxx/4MPN2fnSfjG0XGoai2IwYTDsB3LiITM7OG1VqA6ltLqu4b7brfDvsDkTf8KwqcORVuU7HCrxGOMla+Qzm29KX+jOQ0RAiMJYWLKRJmIicNQCG+sVr1IR3zcL24eHb1247iOxVTBLatzaBlH0Moe7I5mporuApAAEbFD7AG6JGm1utjtiiqgOoC5q2JgACI4+K+19cJXHghBAAxwY5m/8/btf/1nv/+733xzRTGe3Q+rBF51ROLcr9+6ufqdb775y394l8Dv74pCU8EfTCAwsLlUvYQvuy8csU9xg/0Q5OTmyc2bJ+cX5/dO7222WwAgIovYKxKa51hbuf2E/fAlYj9sg5Z1h8gik0Na81iLICJzCwWMoCAAYGZmPrj47Mc9T3pAEZEBhZD3sXVCEObElIgYgQmZMDEmxiycmbJQztyWiIAI506SJGYCNyQkJo8INXcvqm1sWlSDQGrZehkcPQBy/Hc/+OEX/83MmDFjxozHYiagZ8yYMePF4BO+93X8tjmom3Sd8Fol3BSCJyc+80W3IEBA1FJKqcRUxnJ6dqam4Y6I4zjWWpty1txKKc2sw/fuDaWUUsbwIO6kV+hPjtbpN94+vjOWu+P2wD4DACIKoxnUqvfunvb9ApG3w07NPBCZkTAc3CECmbixoY0V2jtFXLIa7kFERGjmgMFMqhrhzGxqrShiY6Bhn0zqphDBRKpF3eJwZgAPzS1buvieG0YMQMcIs70XM17biBgJD0aF4QaAQJTSSAfL16uOzIDMk8n1YQLWUklb4ipeYdsPaC4e04qT2fPBp/Lgszr9djWhHfdNd7DsCNwXAJuOhBMZH97mgU0Y7R7t62hJq4D4XBXQzx3XlUeISMiJylCFGCUNw6BWsUZEEDEikIh7mFkEkEjzrdWq4zC4B0siYvBAsy7n0nVg6uZEbQqt7et71Fz41ZFCm8d2KNuhvpKWBO3uh5iegVpKuPeLfrlapZSaNxEipJxy17maq9ZxQE8RnrqcRAgBMZDQzJJIzh3RZhxH5K6WWmuNcCJSMwRoxV0BXr5H53kg4rKHfOBuufrbVasN2Jdj3bNUQACMKISJODFl5o4abYRItMz5G2+8ebJeL1OSiMy4YDwdh7LbhQcuF11iIwyRTNTnRAjDOLpVijBVL9XHyuod8XrZ38uyFTZAC1CzQhiAGFAQD7LPGV9RCMAC4Ru3j//gt7/xn/3JH/VUy/1PwAzdIgysesSw3d3s6Le//tpH330TUfW9u1t1D1SAgIPqFgOvvGp/nbB/AqZAODPfvv3aa6+/9u67737wwfvvvf9+yhkI3Z2YkRiCzdzNkSI8zLyNLoj2zmA2WaO4GYuknHlfNdrMIqKFudX2uWKIYymlXLqKgYermpZwb2Er2A9p9ps0dTN1KS2QIwBDCV0YkkDmEAAhYMYslIRz4sSchJIgEzIBJ5IskjO1kGS0QLTXqqZqahFGhF1OxS0QB7iolEakmozKV/6NP2PGjBlfdcwE9IwZM2a8GPzbf/u//OB//q9rhTPUdP+ig50OG9Pqjm6GAYKURIR4Ij7BGZCSrI7Xqo1fDsmplgqTU0SYKiKmnCHC3GqpjZ8MD+RMzEi46vJbr9/6+YcbgC3ApBxqRhVq0WYL7pPJZy1azYmZCMLbNCPCYU8cg9ol9RyT+GXaq0cr7wcATVkDABQBSMQI0Myj8WCggUAUbu6GAEykhOB7yvbRCDgooCfDwf0sBwIAiBiRgg5s8fQ3AmmuJUBIhElkIlcubS+QiES46YLMrHlKRwDwdMLNnWO//nTIKX9/b9RxxU0VAfcprthmzNOUbKqIFjjRznsvVmwFDA/cNgBAa4/WIAfDEpv46KYin44SL4ce7GoI4YBJid5+cM4xAABERC11HLayPur7PnddeOTlilgmhxYWYSDiWmsppdaaU+q6joUDMaWUUrLw1lyqOgwDMSOA1qKmj1F6PvIMv2K4UnzylUJEmFuXU06ZTcCLqiIRE/Z9t1wud7uduzFz7jrJ3XjnHoZnYSEs45i6LqUE7m62WCxaJ8bCRNyYFwAARCZu3E3KSQbzvan9Z8beruclxVXS6mFMDkp7pTMiUPNyQiAEJhQ8ENCUmTLRUdet+n7VLwVxmdLrx0cJIcouqgYxdhnLyKUAINdCwFAVTJ1YVZk5PISFERkZWbLIUAq6pfAeYS3MKRNiuGtVRKp7uyQFvIwZzni58LgIX7QYqUDcPl7+5ps3/5M/+d4ffPeb27sfXowXdXcO7u4WrgjuHuqBqU8Bv/Ptt09OTr7zycWP3nn3Vx+ffXI+aqAhBtCDR/71wiXtLiKr1WqxXLLwdrcbhsHVIgEGegR4gHsLvkdEc4HmyQ4Dm1AgAmhfHISlGUyHmdkVeUHL0GKmg5MY7octrYZHy2ObSoNcRrEuR0oEQAgCAKqBwRBEhNQKbu9zwhBbThc2LTYAQUCAgVfwWqkWHoYRwMNNaxUWEYkI3HuLMyApAP3/7L3LjiRJliV27r0iompm7h6PfFZWVdZr6tHV09U96Gqye9iLGQ6HS64I/gJ/gQsu6gv4AbMnQICzJAFuSBAECLCbaC4ITM/0sLswPdWV1fmqiHB3M1MVkXsvFyJq7vHIrMiqyIqMHD0IePjDzFRN1FRV5Nxzz5E4jhSHbDB1P1Adym/z8KxYsWLFiqexEtArVqxY8dKQK2I85hwur/fnCflYapndoaWSIwaJEoTZzIhJWMTBzJIiiTQKmEUkxkWTi5wLHCGGJlSRmENNtaq7OYJT4hjOtuPbb7x2tv2IGim6LBLaIqURx6qN1hkPxwlsEqIEISJzM8cpvoZosXheMtO7mwdRz2e3ntTXwgaBG/FvW6q0LwCEmeDmVmsxZSaqpTr0WUzqE8po8pNLcqOV0e1HmurH+ZQj2BPegwgTgcjchCnFSF3m3L80IXYjR7Q1+DOHELofRmsZ9RPhvjSfLvt0MuW4RUWfTBWfUBveUN5dptt9QADz9qKLBhHu1rXUcGI2r35KrGdmZren2Zhfj4j+NIrqBYGIIczENIzjfHldS97uNtvNAIBIQwillEQkzMJCxHDHMDoTiGKMKaXD8UginIbKdLjeX19djTEw0TzPZlarlpzNdBxTTPVWAWLFqwFq0XZwrbXOs5idn5199OGHjx5dssSLO/cuLy9VlZjrXKer/XSchmGg7aaWepzn68vrBw8eXF1fq/k8z8RsgJqbGwuHFOOQ0pAcfjgeN+OoqubGT+azfinxjBO8887uTRBJBIITKBAz0Yl9TkyBKAhtYxpjGEO8s9lebHZnu21wJOLzGGye5uOh5OISiCElB63MEs1EEcyqmTlMlQCYBpYg4gAzd9G6K2tN5jvmodVTVedcyHx2uGuzEVHcVORWfJHwtKS+e1ERPJDvhL/62sUf/u43//CH3/rqa+fXH/2iHK+tzASoVtUShN29qMZxl4btu2/d+8pbb3zj63lIEKF5/mhffbaeSbjUTV7RT8FvuNudco0xXlxcjOPgjsPhMM/5ZCoGh2nTGMANSyIvWQ9ypqU1rLuKOZyJQeTm6naq8bdpHreukzahMW81b9M2lbPWJ3arNO9Lxfk02+n+G+RObgK0VjlePMaMYQ61ZqdhMKtCVTgwEQzQFKQIMcOstiJ8jDHFtCSXtH2Hw+MQ03YLkWmuWl03l1TSbzbaK1asWLHiN8VKQK9YsWLFS0MdMV1udttMTJvtmc4TnGMQH93N4OZqRc1MyVgZrE130pNnmvUzB2m8iYhwCE1BRBKGELbnZ+4wtVqtVCsFErf3lN9587U7ZxtpwhRf1hVEItIcnw+Hw5tvvvXWm28N4y7nYkBrxnQ3MAFubla12VK3vL6WdkhEEiRIIJKqWkthZjPLJbf1Ra3q7kQIIRLB3KdpcrMY4zAmIjoeDvM0zdNU5qxcYbRYV5xAJ6He6Sfv4X+LnqctqURAwgQI96RGEIOFu6qYnYlgZmTdUhlETUVtZidSmFkAaK3Narn1qy60O3CzwGr701Z3TIu8qJlz9JxDLOFfj9M//UG3ft1Xj7dWp26mpi7SDVmZmqE21+a6rW4t7P7JJ94aNzzHctef+uZpI5Tn5HLpqW/QawYOd3L3Ms0bonHYzKXkw55hMcbLy6tpmt544w2/uir7/eH6Gg6YYp54SXXcbrfHR4+uHl3KZjPeuRBmMydmCWJmQrzdbDbbjURRr2GMIQqtFPQrhVaOgohwpBjZFO7CMo6bIKKqF3cu3vu5llpLqSIDKBp4KkXVtsOYrYbNQEHy8UjMYJ7zfJhKUYBpmo/qCqZaqqmKCIDek/5K01nPi8doWwKYmUCABUZkbj0K5AiMwByDBEIAIiMRbYK8fufiztn5xXa3iUMkhtZ5f9CSNSc2i1qtFmFKTIFghBh5TCEFsZJyhnqzynGtheEMzzkLOQiBWBwoWWpJpqOQD0nNj/NM6oEIMBQASoYKnHxwn2pueIGHkJ7joufAKsgG0KjGNvi8+GWh9eUwPDG9eZF+593X/vQPvrfBcf/hQ5sPkV02KQTRWkuWFIOIgAUsIFG4eh128qc/+u52SPvr6/cezDqpuYECFh10p1E760m3bnn++De/Yu/xwoTVn8cWb15z6bVwd8QY796/H2PKOV9fX8/TDIeqk7sbm1YHiGWZhjiR+xKwHESahFm1LD1nzCzE4s2YQxXMuKmst/1wOLg63OxkysF8e77Q+uuWeVCvwxPxENNAMREH954b4ubwaq7uxYyLChFUNc9BKAUeUohCQUgABtnSh5dCGlJMQxpSCjGKCKAEY6bNbpt2Z9fHyQFxJt+WeHjucV6xYsWKFZ8LVgJ6xYoVK14aKgu+CfqAA/Fms7N58ppikO6oYVVLNbWlWbx5d3q12hohmXvXYq0VAHUGAa6WaylaRUKzoTDAwcQgWBS6c77dDjEyZutuoK3Nuq1mzGzOcynF3VOMVT3PM7M6WdVCzaHavZZaaw0iJAR3atFU7m5WvRKZqqpWQFrAuvW1R3/vLRLLTH2JUlQ1IrRWUCeQMDE9S9X7FHqqDoOZmIgZN7YbCwvcPKB98Upu4mS6lfBHT76kNhPDPvLui+THYLfdRp5QNreXWbTYywp4GQD0x5zo5lu4+Q3dpkr7y3hz+PA21CAICwdiMmoCpEpdyuT0LPYZz7cSfvb4vmg1tAOotU45O0staqXUUkvJVjI2G60VIUgIIAjxdtycXVxgGFBqznOe5yCcQjSzIBxZ2DHEBLM8z6XUYbcBUGod3DgKp1D1WGu1Z/frfxlcOL6scHIwSQgkAlNTizEOZmkYYozTdAwh1FKdKA5jjOl6nmvVYRi3Z+dn53eOx/2wHVnCOG5CSDkXCXHcbFUX1xIiCSHE6O4xxGGQF8Javlr09ank1a6PkSkxEznDBUgSonBkDCybGM434/k4nI/j3bOzIQR2inDUUvMcaiGzwYzgClQ3gQ8hxCCmHIO0LnthCiIM6VVCopBCEHFTJThcQoghCEsUHo2ZSYOUIR7GlNRnMFTdjOAZRo5i7g77fId9vUR8JtyuYhLgxCCAzM/H+ObF5ve/8853vvam1OM8XR3LBKtBJISgKgDArOYGYyer2kIPHMTgsxjffePiD77/zfNfPPjZB5e/eLjX1it0q0bdGp1OBeHl6yt0Rn46HnsvJ+ewmNL9+/ckyOFwePDgwXGeOUQQE3EQMmIQJIYWZ90mSr3/jZrbhjoAW6ZF3BILl20QdzueW0Q5gcDdHAPoKgEitlsRp+1Le0SvCTgCKJLQMinqkZI3WQ0ON3hld3ZjN7AQsbCEIClQCBwDh8BdysA8jMM4DjGGEAILu1UmxChxHCWGeW/FEeKRiP+7/+mvP8cjs2LFihUrngMrAb1ixYoVLw93sXtoSciAEONmu0UREWbyxipqUjcTkTY/JyZzL9pIW6Czk15rVTP35tzs5FxyrrXCISGIRFOYEZzahH8zxCFKYLBDge79RzBTdzdDzuV4PB6Ph2qU83x1dT2kBELOM0lP2qulaNXNMIYgRNyWfUsWjcNbRJ6FIAB0ac9klu5dUaqp1lodTkRm3ijvnHPVqqo9XdCelx8kJtzwzdRtL/oSqC213N0c5EYntp2JXKjJhr05CLdWU1gzdKamZobDXc3MjRRoDtdLZGCrB/jjS8NTW2sL5ml2Izeq6Fsk87Jc7ppn6qGDi/3zjQd0Z8Mbn95drDvrfpKB943fiKRwayvPGrYTRTHsAAAgAElEQVTnW5m/+NV7VZ1zQUiWrZRSajG19qGNIXAIORcRhmMchu1uh5RgXrWZUtp+f91U6uRO5lFC48FqKcm91qq1mjuJUAw5z6X0ss2nvruVZvrCwUxVK5mRubObm7ZOC5FpmpgoxhhE1Jp4zkQkxCQShYNwSGkkr6VUU6+qYI4xucPMSi1VNYjEEHLOpRbgRcjkWz1sKVC9CqDFcANCFJmSEIEEHom2KY4iiXyT4sV2+/qdi/tnZ3e22zHGMs/7y2uq1Wr1UoJ5ZB6YCKiMyUzQjKRYhYMIdx8hE6HAofW2BOZxGIQ557m54ocYQoxBJMVQ3RgwIQ0ypTg4zaCSZ9NKYBCg5kR1sTn6MhGNrzIW74V2byNvrr5jkHdev/PDb7z9J3/wg6/cGcrhIeoEKwDUHeZeLcYYU1BtN1g0AzGi5qPlgfidN+7uLu6+8bMPLn76i/Jvf3Z1zJOqtYCEZZPP4qDxZf1otLN3HIf7r90TkcNhf3n5qJQSh6FbWLG4OwunIUzTnJFjlNbHpWYABWFSAqkzQGjNcA5yQzPFcEFzgj/V7/umgTY1OplAw0F284DTNbDZtQsowAOIncxMzdGqwqcSPgHu5ApTg0VGjNLdkoY0RkmRgmBIshli2wNmDMMwjoNI8/MnNwpM2zGZhGrIBlXf7fT//XcPfysHZMWKFStWfBpWAnrFihUrXhr+6T/9yV/8y/+2WnCr0+FQj4c675uxHbmzUGBhop74xxxCaMyGNPFzF7/QMIxAy+yyxv/mnPOcc55L0ZJrKWpqMIox1qzT8cprllOnLLl77f4Q7oCXXKdp3u8PudrDR1cff/xg2IwxRWF2mLlpXxaSqbmjlMoiLEJEvuxDc4puHtDuXrS6e5CARU7cXBiYW8xVAeDmpVazqqaq5iCw9LXkM9ussfC+5lYrgZwJRmBuqmFqts2LnIcc5LcsmnFaUzUpNC+Mr5+EzUzE0mwP6bSccrfuM03dM/FEfi+vTAsD3Qw4iIl90VnfYpfR9qq5cd/YaxO5dcvn5W26e1/gAc0bui/vTVVrrbVa1RY93/IeG//++CL86RX4C1+TP83fPYPRu9kqt+ElAgkzxRRjHMbRzA/XV0lkniZ1N1WoQkQkeAgAHjx4IO7TNB33+zAOi4+kgCjnXKtKCN0Xm0nVAH9adP6s/Vo56C8K2pGwXGY6cp4jAMhxmqZpLqXUWtvXcdwE4Xy8yvkQo3hhszrP+XCY3MiNj1PGw4cXd+/VUkxVS2GmWmqec87ZQwQwz/P19X6q8Tf3gO4WM6+I6nIpcoGJAyEwonAUDvAIHpjvDunedry7297Zne3GITGjlOnBLyuxqVmpwZ1Vbc5wVObMiMItNrDFkXmrf5KbqblrVQeELM+zm7kqD4MQlVxEOITogKrmnAlox8OBAuOck0iM6cBQYRamqgAMDoc67JYdx4qXilvmS70/yLfj8N2vv/nP/+TH//wf/+FX7p2NXPV4CcuNgiQiZoZ7iCmltLRGmWmFO5hAAhYncQ5G4R8r/+uf/vx//l//z//7X/30b/7uwyazvp0fugQkOPxkEo1X4Yz8DGizGxCGIZ1fnL/5xptEdDxOTGG73TlkESWLuTNRiELEMQY+2V6YgSgEaZXdHnzM1HMXQK27LsTQJ4dPFXFb/Idam4NUK/rpQ9zK5b2OqLeq8ujtaMwUmpEbIwqGIEOgFGSMHAMFoRQ5pRBT6PMshggcau6uALm35jUtHrUELYbq9JP/8S//yQ/f+JwOxIoVK1aseH6sBPSKFStWvEzYPNtG6xyvr/eYpzLtc55dq5szI0po9nyNGAshgNncQgjSG5oJxCEGIu6GxQCzcBwCSwqxlFpKtcHN3NWJCVzvnG3v3z27f2d3eHis1fRx0+DmF5FznqajOpsaaOE/md0JTtQ3DXdqhHNLMSSiTpRad5xYImxg5jgRBN5D1GlxnjilFBIzk5w8KrK2Ftu+a88exK49NgfBGY4Wp0jW7Ayd+v+9G7RttIfjuDO1tC0C931rup7TvvVBeUwoyzg5IrbXuWGebyTKnWPuNPAimMYN5X2Lo+rHoNmV9GG8RSA3YRAZLUqjFpmm5uZqpq300JqVQZ9Ifn3enNjzsrdESDFsx0HmmdxSShjSYT4QfJ6mq6urmIbz84tyPJjqnMt0OOB4xDAyCxyqGiWUfKxaqmat2cxYZLcZd9vtsZqwbDYbU9tfXd+9U1KMKSUJ8nm+9xUvGI0VZZYggUS8VlVNKbW8q1LKbndWaz0ej7XWEOJ2u/353//7/aMH4+b8zmt0fn7x8MHH+/2x5Hr37uiO8/OL/fXVg49/OQ5jGNL5xXlMaT7MpdaU0tluu59YFzPT/0DQK3QAg4QQCaPwNoaBeRvCWUyvn23vbseLcRwkRJCY5Xmu09ElEEjMA7MBUFuaUNqFcMkVM2sXMnI0yXJz0pcQtFQ1c+sBBoATsYTApu5eSoa7EAmBhNVkw7AgMsRpiAAiCMit8YfM2k2FltaWFS8b1KXPADs2ib/22tkf//73/+j3vvv9b7wTPZPOHs7cFd6jLXxJPyZmkdbsUINIv1ETObH3m6wNUd594+yPfvdbOWc3e++jR8dccct8uvcfAY+bY33J4O5g4mEcz8/P7t67++jRo4cPH07TVKuGKGaNxncRAaE1D506t+Aw9xbFscxRADis2WK0PrauMyBaeqweP79OqcmLwYbjE07ANi0REDm8du8185PrB5g5CAtTYIrCgRGEkiAKxcAxcAocAw8pNItw95ZfTWaaZ2Vp9tPmagKiGEmQpwyww//L/+j7//LP/+pzPRgrVqxYseJ5sBLQK1asWPEy4Zblw0fl7muXl4+CazkcS55cq5t6NWFu3ohmpqos0qTEMcYQgrC0oBiWxoZCRGIIMUYWSRI2aWhtjSIRIDOb5+NhLuP5vW9944Ov/fsPP96/P5X5mYxLrXWec4zDZjOiCYCZfKFYW7Sg1irMAIbUTKBxcpE+EdC6+GCkGHvYucPdiUnVaq2BpRkcEzEzc2vUdjPV45FyLnD9pCXNY2jZ580Mun0TpJNYzbGiKaCtR73TooQOvAifmdGpZDDdPKtbJbaNnKyl2+9v+XNjoaKpNwwzUYvyumF9/STD8lvE861H+GLtsQygL3w2dwrbXFVLLaXMtahVVVXTZZhvdf47+e1Nf9KoPeuXn/ScTxeRfdIK/9myYhaJKVFggFXVzWKIh2lqGfYco2w2fQhbSaRWRobWEGQ7bo6yn81STONuh5T2jz4IEoc0pBQheGBFtW43u81mU3MlgKn3ZT+1z/6sH7+UbMWrhFb+EeaQYuRkxLVqMQsiu8324s6d7e78wYOHIjGE0KNB3VKMOo5DSkTI8xxIzndnQUIppdXtttvt2dnucHUJoORaszLLOG7gDrAqiF5U/tgtf9YvNLpIkskDkIi2Qe4OaZPSvc3mtd3ZW+dn2xBI6+H6+jjPQwgomWuJIkSswCBSW2eJSIgpxSQEqzUEYWbrlv4goDXueAIzhxgLMjmqaRAJMQQJIcYQg7qZainF3ZggwjEGYj4fBkopbDYlZ2FODnOtZraUMI0aB/0qjPp/CHAQXOAReGMXfvC1e//ZH//+d955PV9+dHX9kLwOKfXyacuLqLWUYqYAYoxNfptiECZr9jptZlBrzfN+mpXjD77xJrluIv9v/9e/rrkCvnhx3OzDl0z1/DSIaLPZnJ2fn5+fv//++x9+8OGDBw+qehw2qq7qVe1stw1Bai2lFjWTwO3G6uZECCLW+uf0NOtgMzf1JZ1VY4wt4Pep7fe2MlvwzApQ6ysjgAEyd2+uOTcFKyIKQVIMQghMgUjIA4zNmzZemGKQFGXotWQ3c8BYpJRSS2HhlpNiVZPEIQzM4lpbdsZX71587kdixYoVK1Y8B1YCesWKFSteJvhwxPaiqk9W759txWZyi+NIbnWeyZ0cWgoTBREidkIgJhCqVauN+/TeRQ0WnkBwCjGGEDptzBJDBLO5z/NhVjOMd8+2b79+/9/+7ceXmLUxoo/vWJ7zNM3nF3fO06DW7ZM7MWxqZiGEGKKburmbcQhg8mapAZSWiwhUU4BEmIjdrZQiLE2LmnOe5yzMzdyiUT9mRuREMDUG9tfXTv4ES/sUaYgTb4yTQTITS+iZ7E2P3OThvtDFnTpugYWMRbSMJt5jCSG0xRjo5CzZDRBbn/5joXaLncZiwsEnAXT/SzOhvmkNJnS1Mi3qaj9Rte25jW9efuzUmLODYDDV5rttbuquywh1jtgB6lv8rFzqr+SX6dbXX3dt79CquRQPMl3PrLq4mRgzk8NVURXqbh5DGMYRzDVnAoSFmVOMR5C2FTPT4bi3tiB1CiIpRq3TkFJMaX88hhCYP0n+TM/6cfXiePlopwWBVBVmMYYkcjweq6qptUJYzoWI3FCyXj66EokxJFWbjpNdODO5m2rdxjPrnw9q1bQggbk1jlhruWAWZn+RBPSr0/Zv7sI8pnh/t/n6a6+9ffdOcE+OwSGleilash0ndj87GytTgY8puWO26m7u1hJoTVWrmnstpZQqjYRuRu1urlZhc84iAmIzNau1lFoLMR2naSRK4yAiZlZqbUeqlePILTHFGDZjyvPILINDVWvtKk91VyODL9e9FS8PvQjgAn/zzu4H7775499590ff/dpbqdYH712WzDBYPWptsRPdfwPwUppXkhVuanaroo45z6oGQgwCd6gOMHOnw8N3747hd74Zif/ir372l//u79tk5vGa+smL41W/pD9tf8FEzkxvvfnW229/JYZ0eXX14ccfVVNvaYFExBASNbPiVUtPTlZr86DWyEaO7lfW/wFk5CTUU6Cl+XVUbYJlOvnCdc1Ba25rQRfd9uP2KdinXkQBtJG0ZRmIxV3g0pr4mgeaw1WdyUEkLIwoIQUaUhiiDEGEyd1zrlzryYOsam1GcCKBCIDFGGOITlzNq6pJQBHi+ts4RCtWrFix4ldhJaBXrFix4mXix//1v/jz//6/cZCbSxpEN1rmGJjNqFaowc3chSiwtE7V7lfsgMGsqnfDUV8EnNbMcoWbDpeFWUJrfMxlVhAinW2G1+6eD4GFwA59ypuhlDrPmZlTiu5U1dTMzbV5TbsLc0pRK1mt6hAmEnZ36YRDDwqTWtHaronNzKoG4SACwEXqIhRGt8XolCmRsxALMZPpTUTNLTylVG3KHSfynkX0mIdGXwURc3cb7ORWo6PJT5YYdNufuTHVzCc/aDTLUXrsxbuXCNETrKX7bd/hpe/1Zm9vvQ8sJhxtV+n0yk3S7AZwF1z7Y/t54+hxw5k+vvT7PKiY22T080iGn8Hnmrm27EytyQGnJrNadFLk1axUU/VlbFuUFbylWfJC2RNA7iilaFWAOYYU4zwtg0MUYmo82AsfiBWfH2ghi00N7oE5xnB1Ved5nqdJSyGiWisz11pLUXeCM3NwNKWeq9VpPk7z8Y68BrSk0zrPc845DWOMkVlKLsfDIaXUNmr6iVGVz49Xq3zhPVIVMcR753fevHf/zTsX9XDAlLmWdrWHVi+ZiCMLiCtImHvobU+XXS6BIDOrqnBv+mXunS0MQM2qGTETmgOtqlm7lmk3EnInMnjVOoRBmJtNB8wYnohG5g2zCgvJQcJRJDuqe/tnDuvFwleA9/9Sgggt4I7h97fjP3jn9T/9g+//o+999RtvnOt0NT3cl2kaUjTTeTqqNgIaIoGZmhS6U9IiQYKDzTznuZ3RMXBLEAWRAWbg4ezeIN95585HDx++//EvL6d6rFaXY99u4o/H876ieFoksBTRGXfv3bt39x5AV1fXDx89bDGtqtpNUBy1Vnc3Le0c1RvfbaJm196s0xYFdJ89oRPQTb4AIrce1Gxm3YEa3s45X4BlAvbEzjIgoEHCwCEC7M6NgKYmqQDBTI3Re8/a7bulKDIxvFnKw8yIicj746xNEAKxtOtPkBhTCmlQFgNLtSiZdfO5H6IVK1asWPEcWAnoFStWrHjJcCPAKjFz4JSIpZbqJWvODGqJ5M30ueRaq6rqMI4xBhOptVatAMy7/gQgYdFSyuyyWHOYu3kTpxiFyJuQAp3vkjCTg+mWzXIHVdWc51wyTZRzyaVWdYCabE3VSs55msyslpJzbtaNzVvDHTnnEENKw6nB9tTLCaCZfpZa53kmfoy3ZW6bUBDynJnZnoc37N2kTm5k3IMHXYndm68GkREMJKe4m0XpuAiimwL6pIemUnJjRtqed4NRuJmJNGnerfEiWiiYZc277HZfW/WAx0VOfePM8bj94q03tDS0WiO4O1nucLO+SgcJCwQMxeK9Ye6E5zdC/c25sud8+mMbckCipCH5nMc0oJbSHH6HsUwzEw/jhlPyMqvpYZquLi/vv/5a2Ow4BNTKwmqqpsM4bDZbhDCM4+XHH5sbx+AhNpPseZ63anfu3v37+UYw9Xxvf/XiePlgpjQkFokUK1HOs6DVYqhFX83THFMEkHMh0JtvvP13P33IHM7O7oxnO3fLeVLNcC+5tLO41DJN0/F4GDfbRrXUWi6vLs/Pz2utudic59+Aubz5zHirirwKGuiWMVDMQHz34mI7DKh6/eChH6dknsYQokQRN6uutZZc8lzyoKMTtS4QcxNmDiGGGIIonJlCkBBCEIkhwC0Ng5ppgUiIMQ0p1nxs1/k0DMNmDDE6ULSqW6laSt2MI4vokmTotaIW1OLzEVVjTAPTRmQyL+zFvbirGz1xJV3xW0QLYQjEAo/g771z/4//4bf/yY9/P9TLyw/fq4erPB1rrhKCqeY89QmNNcmyq+o0TdM0CUtKw2a7MyeAmsGOqVbNtWpVA8HMaq2QQWXYI93b+Pe+fvev/+5hvc7Vl5YlguHmHrtc8L8kV/UuZzbajGNKaZqm/fX1fn/onWo6c4hwaGkTDYNVNLGxlv4Sp0Ywoi5e8KVDCwQnhwFovWXLxazppRkt+OOmQe2m9P0M/tlb9wlFkQAmVSYSAqNLoHtt34xDD312N621uMFUAxcYk4N8GIYQAjc+m9sMjYWldYiZE4vENO7OLw61ihat9ex4P8vxczsOK1asWLHiM2AloFesWLHiZUOAGjkQgghvIZcEMLyZVpyMa9XUyUGtVVLVqNZO1AqHpv1QUwKJhEy5lOKNLnVrD2NiZnZHmach8b2L7dmGU8CsaB2wtwz+XFXnOR8Px1JqzvP+OJshxqS9bRbNPQPd8VlpcUwG4O7VlKvOpbYHqCp3orlToxJEVUupjdX1pjskLMpWIyZzEAuIAWt/PTlYPIWFyz1xQI1vJ+r62cV1Q3FSDvcnkhu6xcXJN2MhkRf13sJR94RGFr6tAl4cpJde0hNTvCx3lyhCX7bQKarevnoiixerj9bZ2kKZWu1g6SNuY6NV1aw23xIR+IlNdze/sWI82UEvr45nrg1fCkytlMpBylRRStWqWi8P10OMIDgTxiQ2SBSf1LyGGMEcQgBac7ZO82HOU9XKbtN8LLXkUubj0edcSz3sDxxCrRV5VoRqTUv9/HglSIpXS2v72WAt7y5nCgSg1Mru2+3u4k68uHu3FSHGYdSqTJRimqajhGimIA8xmisL7c6248Z3Z5vAVMoco7z55htWsrpP03EsZbvdfvvb3waw2WzkcOR2Kv2ap8izj0VrLv81R+G3hep+zPnjXz44g/Mw5OMkVUVC5BBZGBDm5rDkgLZ7wNJA0qwyThf6ngbIbGbH41G1AE4ENc+1zqUGETplpTbTWEfr0WnPVbe5ZDVl41priEGYUwwphkE4AAkgCRfDUFnqXOo8z7OLPVexcsXnCnKw+VffuPeDb77zw3ff+NZb9y4/fC/vP56uHlg+kjkTvBWhYwAHknBai4o7wkBxTDGFGEOIEoKwNDcON6taDe4gEXGHqoKDS6ySXn+HvvFt++7Hh//vZ+//5d/87eVRj8WsGW/wE87Qz97xp775osMdIch2tzm/uBCR999/f3/YEyGlBAggxGwOIudW9/bYJhOSbpb/bf7RB9nM3U59RScF9E3uhfd05O5CZk4wwM3d1MwUZk/flLz3jbG0WaI7zJ1hgJMzyNzb7IlZ1K0Uc0UgQEiYxN3dSViEQuAYo0j3HqE+YXJiZ2EiCoSYQkhCTApXRnSfN8fhuCqgV6xYseILgZWAXrFixYqXDGHRM2UdzcFplDiIMJtQNFiFKYBaVWt1AgkJMZgMVrV6MywWYRYiZu1+FyGE1qlqpuToXtDMTFTd8zQlGe+eb+6fp1+MfLU3JnoiXMZMc8n7w2EYBjM9Ho9qvvEepE5E7hXdCAIAARUAE1vr5yS4GmqhRYIN7cYRjRZlM3dXM4CaYKd1dDJz6+ElwBw33ZkA8EkJU7eUhn7ietp2CKcMLAcR2cm7ontWGJmCugV0+6MvnbvUfEBIT8Rxj+ixk1EsnWIIiZsZRlfz9HfdZVjt8d78i/HYWq43jC8C586U30QR3lDJTe5kZlq1LmtFR99kPxJsqqQATjGGTw3XF4KDVrNq7sNmozvXjPmYAcBjCnXKNWfPcz0c8zSJhO121yTt11eXdZ6343h5+SimJCHADLUCHGIctts0jqUUERnHTZBIHGS3s4/3bp/dDfuLjlN14cv2xrCIFd1hahUVQIhBWKZp1sMU0nZ3diEiWs2t0StW8hxEHuwP1/uDcby4ON9ttoery+Ph2s1LrecXZ1rz1cOHV1ePducX42bcbDda6scff0xEb24vQow9yepFYrnUfLF9ic39kOf3f/nxDp7OzjQXAUsUkcDEsEoOYhYREDWvDJZT+gAxty4UU1WHgYhYzPx4PNRSW5uLuWWtuZakYmbce/ldzdTczFiEmFq5r2rz3rBaawgiwoGl/YtEShyCZKLMMoEOqqEU6Z62L/zq9iU8v1442hgxEJguNsP3vvH2f/onv/f1e2eDlUcfvjcfLst8hFmKYQhBa+UQx925xN7ehaVEXEottYzDKCLuFmMUEe8cp2njPkOIMRGx1goiZwYHk1g5Xk729t/8Lez4N+89fP/hcarP76jzyh1lBzyleH5+fufOHWJ+7xfvXV9fE3OMkSiAxJ3MnRnc6+MotZpqjLIQytaaSoIIM7dIBYf3uAsnbR7QjxHQ7t0CqxPQ7qZqlWozwSF6xpA70Jr5qNfc+9SnTeha0U+IQGSu1QEHCQViEPeOuSgxSIocYrtGd1FCiwxhbm4/xIwQGQSFFqsA5mEjZfrJ//5nv7UDs2LFihUrPgUrAb1ixYoVLxkcMNZhJipaNuMwbnasE1mGGozdFIBRgZubcYhDjM0Xlc3dnNAkutQEs82cQURiDO7u3q7zjRlQc6tF81woyS7xV986//uH+1/ur1s2DT9uNOjmx8NhHId79+9X83kuIYQQBICIqKqqNVlc1ZZRD2Y2cydXt0a/NrvnJbKmGTQTLfSoL+4T3dixs8ZtMer+SZHqT+Kk7W1uyLz8WwjyZWnZI3ducdoMEQq32WcA5p0xYhZiMnNm6tLsTvjdGDr4aRHXpczUxUY3lhs9A5FAzk43SvD23peu1ZM0+kTTLw9o6Wltg81fNZdiWt0UC2vfnBJFGGhidm8Ls1tNsU+M2DN5/OcZ56ef9SuX7s94gDAHEajGGGo3DQcx3H2eJnNCraa11totSISgNedZS9YY5nkO3MRQomqHwyGlNKRBREou03R0M7QPlbupNjvt53tHX3B8oXnMF4ilqwBEAFOQEGO4fHRZq5WcTbXpZ4U5hEDsWrOqNjWtaiWieZ6m45TnPM3zRZNUlzLPk5mlmESkXTNLrUNK7m66lOE+A4v5iZ//U1/60oHwheagHchmD+e8z7mU4qpKXlVr1WymZZ5zDjGICN1EkFHLUCUgihAHNOdZN4eHGISo8Ya0eO+7N/N3q6U6CCQGqFprX+AYJUZmTrWmlCQ0VaY3m+qcc4rRVBmIzJGZi3qtXpXcmYicGJ2/tmaf/wLOli+PY8NvDL+56S1G27dlwwQIcDEOf/jDd//kD/7Bj77/jR2U83R3+ArhbWaOUVIIQVhVQZAQ4jDEFEMI7Y5oajnnkvNms5Egaq5azBTNQMK8moOZJYQYAZScVdXhJFLN5urDxfCPvv+tt998/X/5P/78//nLn37wYC7m6k+cebdK2q/q5bTv+TCMr92/f3F+7mY///nPLy+vTd1Dd10z62GtgLcOuOa8DoSTFMBwU+3Wm4q4wwm+nOnAUuRGi/NtE57AbH2ih+XPzZT5GZAgMQaYuYGJmrk8uzvYW8MYgYjahyTGEAVD4DGGIIhCEpgDkxA3JQVx453bbSIEDjEQwVzV1GspR5pqnSuCX2X7pAjiFStWrFjx28ZKQK9YsWLFS0ayUAhw2085hdJCY7hRnURgbssIg7MIi4DZ3Y0AYREWsLWWxiYSar4N6D2SjdTkxR+DDMI+SnDh88Rv3T2/s3tIuF7UwrdBrYH6rt+9uDhn5nkuZnB3EESkllpqbUx0znlhekmbFTWzmqoqc8tCpBML06lYnJJvQCAWVlVzBdBz2LtE2I7EGVMttbfR0omMvW3Ue7K+WAjoJjReLDXaRpnAJ/8NAoGEKDAz0+3wQV8cOhrboqonC47T4LQvNzplnLhkOr2FhYNG109zF1L33ffFPNFPe0o3y+ET/dyWWf1FUd1RYao9kQdOIDc3dmYyY7oVB/Ti+K7Pg4IhAjyXYjnnWU1DCFoXbxPun/yFgddG2scQBAhBmNhchSXEqF01TzXPZZoIKHPJU06jws3y3JOUvgxE0jP17F9ONNZDmCUEY3FUERERImHmpRWDUxpijK1RwKqmGGNKaRhE5Pp6fzgcVVFKTSmpap5nd08xhRDg3ixox2HYbDbMXOpsn+2c+VLJK9V9X/VyzpdpHs3HwCRCzItPhhMhxMgsN+9niWMVJgnsoFJKj6iNA8O1ZAKW1nvA0aqYzMTCxHnMEgQAACAASURBVNSKdMztZsZEZGjbai07zIs3Umu4N7PTBbPHprVgNGGFq5sv/KKfLtOn43TrWyzfPnVknhBwvvAj92Jf8Dlf7YXcCfx0byOiliNJS9gBOwLhO1//yo++/83/+Pe/871vvPXWnS2XCdG36c7CEgovZl8OdzgLu3sp2c1hrTrby73toUTu1oyC2YFSFcQsgUUA55RqyaoVULMSTCNb2sWLzf3rH333fEj/6q/f+7uPLj++mrgbQdwMBBGD4K7oTVI3nPTzjdiLPY6f+bLTPuG73fbtr7wtQY7TdNgf4BjSJqXRnWsb434eERGxEIAQQoyB6NZMoQcsO7cbZTuiDjiFphjo4RhwQzs6LdWQACLpUuplQvTE2zmNKoPapaQdYXMnGBFJO8fJA1FiTkFiDClKbLwz93+tvh7kpots+UcgqDu0grzNiNTcvBSFu1/uVZ5ZfV6xYsWKFS8DKwG9YsWKFS8Z//C/+smf/Q8/SQMOWeX6OJJZVbZKrs05uOWtmXtMgYjUtHn8ghEkBArTNLVwvzYfd6DU2hYNTMRETkwEESFgCCwcXUJVf+vu+cV2c2JB2wJi2S83t2mazWy73W63u5Lr8TipmcPbCqSU0pigaeIQAnc5jIMQY6pacy5Njp2G1I2MTwxs79c2VRMJ4zjWWlSrdhVO3yc3Y7A7VA9dr3MiER7noOlkY0Etu5F6BDzaMDSOgkQI/bdgoiaf5GWB1QYNy8+n4MTbbacNBGqynSY0ctxauZ52vvk3uxOImVnkxNd0fvqWapp6Q7r1t/aEPvq0tDOrTRVoJ/ra3Q1m2o7/LXL8cZ3Xr70Go1tfn/lXf/yRWDb6aVsspeyPRwvh4YeXfr2PjnEYa5mGYXj99TfS7sxjmqcsHEKSIQ1wIISz83MtmQnDOE7HfdWqQDrbff3dd3/6b/7NBx984OZ37792dna2v37EROMw2i3D71ccz09SPHEgXkm0YFVhDiyl6WRLOT+/cNAwjO2UFOFhSMJ8PM4sMcSoRSSElBKA3hbAPqS02W4Az/ORmc09l0LEMUQtVVhuiJPPyEA/jlM9rKMzOa3XvLWmf4FF0OaY3R7m/Mvj9DqLM0sIHAK7NRKrXS1FhIh9IXvapdYB4ZZOUAEiCUNKbpqPBwYFZgbBDW4pxdjk56ZEzSKAQwwppXa9rbWq1tNls22OmYOELojuVkvUw3XdnODExa32MAGcinkEGLhfB8keOzrLN/wYKX1zuTjRVs8yFXgGntvp+0Vdjp6ffX4xnzoiJ7gBTBBmVyNyYSLzKHwxxD/+0ff+i//8P/nBt7+yYZsuf2nsiMxpY6qtmlhrMdNm1VVrUdVaa8mzVnX3YRjajbyUHENoktp2FjWTYq0FIJhZabd6dq2aZ/NatbhWrjGFlOLwJ7/7nXdeu3+e5M/+8meHY1b16l4BR3cbIxIQHNa9uJays/UC+KeP2Etkn4HFVAzA2dnZO+981cyvr/el1BDSZhNCGsxcqvXCe5sALsO47P4Tb6FZnFgr+jSjZ/jisNOnba5Fe6OVw0zdXYiJ3c3YXbsK4jGZPJaCEPmNPxo3XQQx3fDLGJiTSGCKQoEpMgUmgjGkJRa2YiRLi4m2fjFteR9VS3UiiBAHYZJjrpVDIapXG0sFK1asWLHii4GVgF6xYsWKl49rXPDDy83O5lLOz0arUy41z0chF24LCEgMzY+vzblbA6K5F6vExE5mHkLobcvdPVizqqqWnBmUYhQhgMzJHVH4W+9+7Ss/u4z0s+zP4BAJzkLunuc8TdM0zfM8q3WKpjERTQjDzAsfJI2uBTywUKKmwSE/qZC7AtnJqrk2M1HUUnJfi9YiIi1rrpaap2xqeLZ9whJ1DyyOFgYnJ4AdxsSyLJw6mu10F9A5WoM/N3vgxRwaToLWbgq4g2Dm1hw2bi3cWhohWvJ6f3lfFmuAU1tskdFJZnRL8bzYaywH8ySJPj2mv2LXSS8ruvYAAgurM0xvPdhbh/tju9N++Wkfvc+Pmf1Vr9zoA3hKSXZbOx6O+ysyPx7205w3wOsAMQFW1UvJVguPWxC5Ggc5OzsnV1XN+/3AVE3VbRjGNA5mNaZIxA6HiGy3LPlZLMyXhpX+or2RF7RLDlUz4DgddZ6hepxqmUrOhSVc3L2n6sfj5IaLO/l+iDUXczscDjzPF/fvxxgvLi7mw/Hq+lBKvb7eD0PMOe/3e3cPIg5XVTM/ThO1hD3hZjH03PgyEP1P4HLOvwDSMIzMI/MuSmBiIndU1ZJzbcbbCy/lcHIjM3KHk6k6OARvCuU8z0JggrfLeymoLo5AzuQOmFkpJc9zzjMHaT4MtWoppWolIJfCQch4yhki0X1SLU6h1uzIjmOplzk/KqV2w4Hb10yg+Qn0VpHPNhSf9fGvPha7qsfeuN/6xkEIzU4F1pN2zTeCb37l/j/70x//+Pe++85ru+ODD475oPPBzUR4HIYlnxeqtZayGUe41zIzcxQOKRWqqgq35j9cpim711qqmjtEQpPhm1tL/G2zjpgi3My16qyaVWuUAHBxUt4k9R98/S2tvo3hpz/76PKYC2DMChQz9woQ3fKouvHq+mKfy7TMQ4R5t92+fv/+nPOjBw+uLq/3x6mo2X5qD6Q+aVAW6a7NqmZOt3zJcHoo0AhoZm5x1q37wW+Vw63WpkVWrdYiKJpewMxMe5Z0mzg9LoIWIIqkECMb6yIkwKIRAMihVUupFCWgd0gIKLCkFFOSGFiEQK61OtlJAc3cp08tsTKEAI48jhk5G9zL9j4dfhl/C8dlxYoVK1Y8D1YCesWKFStePo51OOx++K7/lTO2u+1Uj5oPLY6v22cwE6C1mvmyJEBT3wJNqEsOJem9lu5w01KrA6qdpmyPbk3MFClKuHf3/O6d3XbkKXtRRydmccPWueecr66ujsd5mqZ5OjbDDBYWCSJySrpjat3SZKrurmrU9MKNDHBf2OdmfUHmXlVLruZGRLWqqVWtqhpCaDrgkkues+rt1SA9pjO7rb49ka/U2AdDS2jvKxVucqcmbmprHhZu+mVgsZoFmvCZTrsK+CIMX2TSzaMZ5k59tBcivP8RfupuXVys3dElyu2HLn72W0PSGO9lrPp7unHKRtdbO1rY48nK4wadbl7+0CgXpycfdnswXx46gcXDMLANWjJCMNh+v1dzCQHMcGdia5bW7jDTqmYGFwJKKY2zMC1XV1cppd1uF2NS1RjiMIwiweEswXsf8RObX/HFBbUTl5lYoNSZrxAKyjAMMaZS1R2qpkUJFGOa5weXl4+IfNwM03wE3cl5nqe5llqrNivhEMIwDAeiUkogGdKg1WJMqgYQk3TH4V+fgHr25+oV+rQda30AXBBtOZzF7u7fr2cG7f04Vs3IGS0Fl6j5upqTWUs+cyZSR62VpD2M4VB15nb7aqpwJmZzr+3S33WyaPLIZjCt7sWMHMVcHBnIxJMZFd2rXtX6y5yvSp2rmfcLsEF7uw0WieSTh4CWy+SpEHhDPn5qVeEVOpKfFe0W2Btolnfut76ik/nL7wQYIp9twnfeeeP3vvvuH/3w3XfubyRfHa4e6nxAzQBYpE6xmUC4ea3VTAWuVo/765RSECEQkxvMW7MR0EIpVbU2W/YY249YaGIzYybXRESAaZ1LnWrNxuJgNShN4vH1s/i9r95NZFLr3314+fH1VMiLw/on62R6dSrWfvLd8guD9hFk4t12e3F+vtvuHv3i7x/88sH11fVUVPvMhJm56xDMRISZALRkz5uOsQXtr2ZdAW2qRMTCuBWW7GZu2oKiVRVwIm5tDf3q0IIBn7qANgJaAO6NY2ZmcCOCEznYfekngxOaIwd1752W4aDgJi8QAAoHSZNhtNwLJ0KMoRHQSswhGIoRuHId7F/8xV/8lo7NihUrVqz4VVgJ6BUrVqx4+TikN97GzzmEwHJ2doZyIJ02Q4Jr41WZiUB5nmupjQFQVTcnYpEgIbA4KTfrzDSOLW2mlFJyLhJ43MJdzWotWmtRTTGGIMFpM/L5nXD5oJI6tecvbeLuXkvZX19/9NHH7si5HPZ7EgkxpWEoNddaAbSVYYyRiGqtcCdm6VZ9neE1s8VGuf9nTktIzuItoT3ORqQwzwBMteay7E1X/bg9cwgfRyeA4Wh0hrTe4RaC5csiVtSV1Ny6AmdZNZ0sE5sC+v9n702aJLnSa7Fvuu4eETlUVqGqAFRhBnoC0Gx2N0nR+AYzPmkjM235F/QzRJlJC621extt9UzSRqadzGSU6Wl4MkrkI5tNdpONHjA0UGNmxuR+7zdocT0iM1FV6AK6gM5uxQEMyIyM8PDZ7z3f+c7BrUNzfXUMwaHNV8VohkgbFw+ATcLiViZYwxdj+5G6RYF1fwPRpkn8HAFd+eaq295Q0KNxdrUIcdxKni9It8Yp9SgR/9R0evtmfOT1x+ILi8Ieo6k/v1BCZCYQ3mwLQaA7VLkkOoRq7gc3A+K64b5ahxlt9jQTN02bus5FhjyM+vXwCMg517pD5RNJhIh+h8ijz7Uh+Lhj8aWSLHh2Dv76CAeE8HDVRJhEqrFGVd010hChaTXvsSTiYNXI3bSslqu+XwNQ23aAVN0eqjuHuRVVVQPAlBpVhajFPvqVa/TkrX7CH7alj/EWdqkZLo1Ym93PZb+x60RBGAga5gEBiMgRqBZDUSBKACLMgeZGNfYU0B3co1of1dC4lKRtW6J1BJIkkaZJKdyJOKVENHpguLu5EWFKqWu7lJoIcMDiAIQuyZgzUmHpTUsuD7PezeWjfnBAIKqnCmLlMmG7u0dOOc6OEALVO34V8Qaena64aSTZvvURNfDvzG3kPLbs85O2LsYHIoRZjJQiwtWpvP7C3n/8p9/7vW+8HnkxPPgoa8ZwcAOr4YF+ala9vtWUiJOI5d5Ml8tF13VN2yYRdw+zGO3FqkqXRBITEVGTkodbNYMOwADVEgCMDgEehmGupQyDIjAl5ka1Dx/E6dZBe9jenAn8zT/i3/xTv3JzgIRg20L++LQdRwCX+uI8BxE5Ojo6PDwUkfli/vDhw+VyYUHIQiwsjEQ5m3sA4DbNOQAACGDsTDtb3DjooMoSbxHV45sgPACRsDaIjF5nIgLuEG5uY0CIf3p8Nhb7631BzdXNfMxPrpVkZCACBBGShkXqkJZFiDDM1XrDIZggNaMaWoSIkZlEOKUEEIBeneUBIyKy6eDuECfs+3knf95hhx12uETYEdA77LDDDr95/Nmf/dn/+9/9l26MbWS11Ex4msGKm0YYbTS5hFi4xIaF3OYtlVLqK4QYCOZGo1keVzsLdHDVnDOEI2HCJrUdNo1Dc/3alVduPX/S310N683U68IUtOSyXC5m072maXLOgMTMKSU0q32a27cjIgtvOjJHLduZ+8Q5IgYRt1ad9T0+2loDU50djaphRHw6uqYqiQmg+h0SIZIkYkIABN7Mp2DLL2FV8mz4hoAzqleYKw9V+fEtP0JY318D4TfBgBF+1o8+zt2oxkFuGe3Nn+oHMLbuIRvJ9Bilg5U1x0qLRG0RHkXfG4OOoDOpNDzOVmIrXXvsjntK9uTZvu3TCABEYhFkMfNQNbMIjEDhZFo0a5SS+8HMsGZRAeTVyk2rNLL6O08n0zSZDIJeW7tVPZyQhqGvFZpwR3cWwZGA/urJo0fEl18cn1EzeMpywleGx67P598PG1OaUf8YiYlUzdRqpaxtmgi3cANoJB3s7R8/7Pt+fXDtqubiaggokrquqxeXe5h7RKSUtOh6vXaPCOOxAFRzRy+S9s8I1TzncRYHlw4acaz6sOhCda1G6KXvzU1Ccs5ViOru4YFCiYXcinqgI7KkRIDStCzJVXGkpKOU4m4R4OZmpspWyjCMVUwihAgEYCSPMLV+6HPJgJTNyDyQBiQLzBrzgBP3ufrdob8/5BJBhFzLjAABQEhA9QYcAE4AuOl62ex+D0CvDgwXnzAR50/Tz6qi/S5ic53G9jQ92/AIZwQCiICEMGvk219/9d23br37xgsv3bgyZc02EKo0POmmuR8Wp6cigixM4zChScnN3K3kQd3MfdWv10MPAF7dcMzqA1a1RAQRV/6UuBqLgZmFe43PQ0JmVlOz4qBRHbbUiKRJk2LuQJxaSTzr0mu3n28mh1dvvPB3P/n5h/dPTnO1Eh8v9N8i3nkLZn7uuWuHhweIeHpyenJ6AkQIhEwpSW0yExZgqEEdNYmXWRCx1AjBcwT02Agwtm1BeDh6NTypf0eAsyjpOtgjFmbbdGWdx7YtrIIQGyJBRHcMZ4JGEnjgaCZeg2VBqFLj7qaqQUAgKDXEmoApqokIANWRExETMRJBWESoKQUxCyVxCAcwwxeX+/Nm+BIPww477LDDDp8TOwJ6hx122OFSgCIa6E3bxaKfJEIWt7Ix/YWIMXycRcZ5U+U9kcJDzSC8qnMBwMI5nIGqHzQSVRsONgIQwiBmIAxwYbh2Zf/V2y+89+H8PqwVzk8569QMi+pqtbpyeNR1k5RE1QGxaRtW3ZhRuKlVXpaY6oq5j1mJlXgGpNGXc6MRpsrHIAGCu0fgSBYj1i2FCASikKAAd2Zxr22eT0LtHT4nVGYmYcIaN0hUxctcbalHA2hEIMaoTBfWRlMQFkIcif6xeXyTIwbbf84kyxcIaABAHFtWzyms6kfPpnnnXt+qwgHGqTASxnYRW5a5uoWEA25FlF/SrPnLZZ+3n8YAMiOi1WqFw3B4sGeleXD33jD0jSm2bdu2TWqUEBC566gvZm5ujJCHXAsX4R7BQz/kXNrpdLp/0C8WbdvVmk09TK7bcLLfCJ4hB/2svuI30mn++VYSEYWFU4NBgNg0zZUrV+58fKfvczvL7s4sRZUAUjfZf+66Df39Tz5YrZaUuJTirR5eueLqi9WQ8xDhREm1LJeLCN/f259MJ0Q0DOvjk+Mbz10XYfdCQoBPv5K/gljfsjwX/AwuPTxi5X6i5X4eruokEahHvaPWiNhtXbBmAwKAW4CMtT9CJpYtvVXLfGbqHttdWx2lzdTMsFZYYXRxqrc9Nc9qQJE9MMID1oBgAEXvFXswlIdZj3NeFt3YCwMhjA4OCBBRTYqFsEt07ejw6PCQEUspq+X6/vF82Q/1wPm5rpEYy31n0unNLtl2jfyuMtHxyI/n9OIAAIEQBNAwTZt0/XDvpRtX//j3v/bOm7dfv3XN+3lenerqlCA4CUYKt1JqwZtqsDDAyISq6lCKheVqvGW1JOQeDh7CwpJqtgRzaHHbcNA1+jgiaAwg5AQ4ZC1aiIOFWZgwRNpmMmOPACRuUtumZnJ0fXr9RX7ptTLd6w5/8cuPHqyOF8tV36u6R/jZDfGyX6JbDlhErl9/7vDwQLXM5/PlcsUi9dJjkTp4QEYiYsRSwAwRQUTG4vqFIQSOBTLcVtlpe7tGBETajAfHujYFMRMzu2ls727jKGlUG2w5aEJM1VQrgAGESJiBAgPGaMEaRQhOYwnJx1Y1YGISQRYgDMKouoFahB6/NWoyCkY9kuiEPOSiiB42b9f7w+QrOTI77LDDDjs8FXYE9A477LDDpYCAFiQr+vHde9cOZzQs82oephgGAKOQuVKUETXKXM2YgUUms2lNma8emu5eTN09pQSIgGCmBkaJkNEjAmG9Xg3qPD3cnzSv3rp52P1cAAw2wtsRCACmmvs8m05v3LxBzPP5fN2vA9Dc3FtmdvNSsrsjoqSUUiKknIdSVE3Do3q5VgKCEIkYCX1smvdAjHA1qxtVyhhCOJqxNgCBKgLh/eCl6JNYrNgkotcO06qGoggiIgwiiFFjjG6OhEBU1y1G3VxAVdIx1biecKfK4MPIE9ev3gQp1gbVM5J486ZxBrbRK4888paOiY1iaGs5vfHGRoDRwrl6SVShe11QfQEdPWwr2X4Wc+U4x618tXPvqI4iARCpaawM8/lC89BNp8HcTrrAWPfLIffUtswEEWMlIMLDixYzHUouWtK0vXXr9p0PP7Cch9UqAE5OTnLOnXuYgxYw1ZLN9CvdwEuEx8puv+Ij/rmZu4gwN9cS4UwUpsfHD4np4PBgf2+GiGaqmpOk0JLnp8MwhPtsNuMm9X1/5eBQqoepK4ATQduknBohQSRzBwhm7Lr2uavX+r6fqTFzHnI8kwvr3FY8w6V9ZYiI05w/WC5fPDw4aBruugQ4absmpdoAX9trWJioPqMAiRHJzR3B3bWoqoa7MDdN9VJAImqa1DRNSslKQaTaRy81QYyZiAKDWVJqHFA9ClIgK9AioBQtah8s1/dWq+N+qHT3JCV3VzON0WjA3SKqdwh0iV94bvKn/+L7//yP/6hpmrt37v/Dj977i3/7lz/5+Ye2uSX72M1SzfnxrPFma80RAUCPz8L9ncFZcZc3z4Uz65itQ8dU+K0Xr/yLP3znT//4uzP2GBZ3fvojCrXcn548hHBmTql1Dy3qm3GJqpo7IY/RERgKbhHVmp2QK5tJwti0nBoOEJGum5Zsql5TAUS49kjVjGJmadu275dFhyaNS2i72XS2v79/xQOy2mq5BiKWJjUT5FZD3nzrjZ999MkPf/Kzv/7BD3/8sw/ungxugQBULVkurxg6tuRvNddKSZ5//vm9vdnp6clytVK1pm1ZErJUNwyp/RwAHi7ALMTMABABDaU67NhYrtfeLDjPR9fSeDVPI+I6HqlP7bpC23I7bEvq5/6yKVON+zYRCxADJBKuGxBny6q+W3UbkZGFJHGTUpNIGCsBzRjMSAQiQqM5dKiqWiRhFg4gDy+lOOa1mioVMCP+87/4i6/wMO2www477PArsCOgd9hhhx0uBd75sz//d//mPwf3hZd97ZJHUQstGIpIpZSIEKldjKO/AyIwJ5FEo96XmbkO7N0cwoFw7KdEABp5VYqIiLZtWDwSHUy7m0cH+520BMXBHlmxiDCzMTfP3d20FNUxsjDMEFFEtlPzMAuKJEJIyXnkhQkR26rhBqjWCK5qpSjL6HdR2XOcTkWEmLSoW2VvcSAchp4ybdRpj2IjwgmkqjgMAAsPC3dDRnQCZCF2NHNEIEOPOK+AronqNccRANydibbOzrDpzj7HSI8zsHEVRmuO7ZsD6qaGwzke6oJ3BgJi1X3XmSVW/43xnV6zejaSPvBwVzMbd8sXPdUe2WkbfBmM5BMpGzVdD4OrllLqbqw/rPs1irSTDsMms3a21ymQu2FAatvUJNfRkaZt22bSsQiYBQTWzCWz6vObe47wsIw+YChtTC6/cnx5X3r+eH2xb/nKOOgvsnpRTYFV1bTkAUqezGbZymBDPwxpqsQEaBFgOpRhlRIfHB6cHBdVmzVN0zQPP7mzWJwG0GTSMqGV4qoEwETLxbw7OEzgQ+6HPDAxEtamjM+5XZeTrnoG6N0f5PzJatVGHEBgRNFqf2LqplrU2J3MDM/RWKolkH2MKvSAqnQ2IkLAWiUN99FGB3Erha4VtQB0d3XPZhRRkNaBRaM3vT+UedGl6vEwrFTHBhpAG9Pq1MBHrwAIpkgEt1+8+frLL3zrzVtvv/XaC9dmbds8dzh58ea12Wz2l//+h3/9dz9crEsOYKrVjjPHp4v+BLCJM/xdxafFsAjVDB0h3MEIITFOmuaN2y9867Xbv//1l77xys0Xj2an9345f3h3cXy/ScKETdNWT95aioBzoQhQn4CBzMLCQARMwLSpxI5lWEnCJLVEXQ0WVMMNECk1jYjUOjcRRgAxNakZhrVpbhIJExF5EEvTdBOSNAmYzvY9AJFTaiNIPfb3bhxd2b9x4+pLt5//yfsfv/fBgx/95Gc/f/8jC9jS0M/k4frscW6lJl13eHi4f7APiMcnx0ULMTfEyAJAAV7t2AkJMCgAkQGwpkZv9iEhkplFBDOPJhxngE0f2ehZVmnoR/l5PPepszUdLdTGNi8CoMCaQ4ijAVlEOGDAOGgKQhQiYUzCIpISS6p+IUEEtTYhXDvYqlvPWZCiWqgWNQ1ATIwJHBACCJp4zJB2hx122GGH3yR2BPQOO+yww2VBoDpzOAYiihCiQbgHUaiqqtbkd/fIOUe4iAi7qTFzlR4zU03oKlq8OnWaOQQw4dhaCeERZpOuA4ABeQ/k+uHe0ayZNrTq3R8hVKryJee8Xq8jfLVcrVbrnDMREXO4i0jTtriJPYzwOl3EjZYXAAAwSUqSmMXd1LQGtQNgquHlzOt1r6pd11aefaCsVjloMDNiGgmLx0wPH6HhRpo6wsDHpk4EAHYiwahbWSoFXBnr2iBcp1y4NUPc7M4tJR1bAho2zs6VQT6fUngmdga44KFRRTsXpmqI6FspNADEOZ60EtAb65LR7UNV1WzUUG81UV8Ej/3gsyXUPovLc3dVdQB3x006HIaXkhGJmTEiNSxCpZiWEu7UtsiCZoQIASxCSOEOZvXEY2ZpEhK3bbNAIEJhBC8MlpiYH5sv9ytcFC43Pi9b+qQXny3h8mwsR2rVDEXQESAIQEjC1xYQ4TVwsm0bjFojK4hQtJRSkKntOgDIJasWJDEtjXCY5r53tSalIQ+mZVNfs+lkQkhmebxYP8f+ePSS+S09lz6N4j5X/eVi2bk3bXI3Bthw0FpK0STuaXP9IhE6oJkFgW9SzxBRzVSrk3sNtlVrHDa7ySNUrajWm51FFPdebaUWHhlhEbAuuvC4ux4e9OvTnB2CkBMnrB83Mx8d3wGAENrEsy5d2eu+9+6b3/v2N37vm290AqFrcrt+dPT6qy9du/7ctRtHy/70Zx/cuX+6RAyLqn5F2PgbbcSmcO6X32GcP4cRiRm5GmUTxt5scuVgeuNo9iff+/Y///63v/O1Vxof5nc/Wi/n/WqBEJJS27azvf2u69q2dQgkpiRJxoe7iBCSRyAg1oCKJJwEiWFTfq5jiYgwc0kcgKZmjhBUxc4pJTMb27zCq0VPyYNbaRIIMwbMFys11zwIgKSmnU6rSxMRl1Kg5G46GsFALAAAIABJREFUu3m0d3i4/9LLt7/xYPGDf/xgyOUXH/xyNNn6tR6pXzLOuYRMZ9Nr165Op9Oievf+vSHnulfNwcM21l9jiAVgjO5hZ8OPMV1wOxTBTfh09UKp+SKIURUDtYBEZ95fZxjHSu5wrsR+YckABMABhEABBONgBmDkwWvVXwiTUEokUqnnMTkYwas1D2+irbWYRxAiBiIBIqhqqbf6pmmkJcdAgmCC8DE1cYcddthhh8uCHQG9ww477HBZgKXniSCm6aSdEqOu88otBzM1TarMZm17VlUzAwiWhMilFHXTwZIIMyORmwdEbcBkAGCuomNXczMrOREQYph1kq4d7r1w4+Dah9P7nywemXyN8+/FasUnp4S47oecS84FiYg9wrNqn3NVK1cVYWwFKmfqJyCmMU6GmQh14xGNMMq3ixZTmy+XzMzElXCPCASsHtN1293UwR+dCD0NRpHdaDToVLnnDW1RCWN33PhqhLuhIlKVC+GWgB438JznxshEn9PlVPb5zD9zI5aOje/EZu9uKXoYQwghxij30YQ6zllHx6grDN988kLaz+dhzp5Epzw9zfLod+HFn/GRP8X2N6xmLEwsYhGE2E0mNgzT6WxQzVqCqRRdr9fZMTyqEM7Cw93NzdQMh6Fvck6JETDcAZElBZG5qyoTt23jsAksqpq+x9OFT9pvz4p0+vU52af5+AUW6Yt+0Vezqk+xFERm4aYVaLBpawcGIjYibduKJDNr2zbMEAPCSykPHx5rznuHB7VTpG3brmuHXFbLJdPmHmjGLMxj7ahpUtsmFgGEamD0hbb3t7qM8UR4xCfr9QThemJw7yBSk4jRPbC23BCJMBGWJEnEgUTEgIgopUTuSVKTkkhyBwBiYmKu1UQH93AIBKAItMDBnIpltT4gM6tFD3qsdlyGk1xO+35tFoCMAojqHqN3cCASE6mXmoVw/dq1d77+2j/7g3def+nG9auzBCURNFORhhGHfv3gxnPTf/Uv/+Cdd7/2b/6H//F//l/+7cOT7B6C4AAO6Egj0YfnS5u/awf3HGoYAoDXCFwSlkTipU8EXdf90R9+57u/961vfe2VN28/f+u5K1O0vDy1/cPX3vqml97KkISJCCMqRWhQwwoANjLYauOcJNUDpgBRFFSJE4swUQRYQF73Q98PQ57Npm3biQhgWJgWhTAzQURTK6VURy9AdC3gquREABGr5SoA26Yb1ovC0radmau5OZSiOZdyNxRQQXqUk1VZrU5zGWwsSgeMXhCXjoRGrDYVo3h4Nptdu3ZVRB7cvfvT93567+7dxWqQpjUL86gbgVsNcqWDIzACkICqh5ejB3DNfHYirrmFYBZuUN/JUm2v3K3mi4B/eujl9c0XEZuRT2X0CZGJBEgAuAqix5Y9EqZE3BAlRmZgxs3tYVRG1zGQOyp6qLOTGbpFcVcb1IuZQTghNE0zmRzMDg5XqmaBEZDgv/6f/q+v5PjssMMOO+zwtNgR0DvssMMOlwXome6e0NVbbgpNg8RE5IhmBgAiEgFuVTlCIggQNVpPhD2oKls8QkYuFKulphMhkYerGqAGAoW7VxFbBLQtyXOH06ODCX2yoFH/FxtytDKhvlgsCLnt2mEYhmEwtaplAhgjY6rsBZHc3cwjnIhqY3s1QqZR7oJEjIg2GhxX/+MqjquEs9epSW0OjQgMcHM1q4GGnzk7jPPyxeqrHIiEBFuKmBGJACMgRivBUYkz5uycdSPH6GyINDLLlTne2m5sJ3hw5shx1sFfTTJGgprOlllpr/MyK9wuYkP+bXb7uEfq7LEKBHHcrI2J4uVyAXgSd/nIiwFC3CYhLYnZAIahN3NQBaLlclGEnifqh8HMum62t7+PhHlxCu41QtPM+uwzCCJEQBEpuZwcHxOApHT88GEppZQyFE1tG1hy0aK6WZlLs8OeFk9Jfv36TOgl2jMeoaX40DNGcS/DwAGE1A95ve73j2A6mT6882GYHlw5SikNfX7+5s2HD+7263Xf98/fuDns789PTizg6tWrw9BPuvZw/2A1X3xy9+MXX7o9mUzcfRgGc18tl7OjG5NJ90V9Wn4bT6pfjYhYlHJ/oDtDc4Qwbev9a+wLgXO3qapLBaLYNM3UvFAzc+fqCBzugDB6JLmrFjMLRDVHteKhxXTIg/nCYgmsRedq9/phXnSp1qtZZTNh+7UeEQFOQEw4afjK4dHzN65/482X3/36q7//jVevHbbTBt36NnHXJk5SWbamw2sHs9vPH9398F3My5/+4u77H97/5O6xQhi41TiE864bAQhn+YRPxvm/fsb58GxaBD4PHltmu6h6xlr5BAJP6J04YTx3dPj6q7f+o3/2B9//7tu3bxztt9KE6XIdWkREmkQwJTCMqG5T9XCEW7X+2vT/jLypQ5ibqo7ZsA5IVr02asUo98Nqter7vuShbdtGUq2w1hYoJg6IelbVGry5gxu4kSthQHjf9+5OxOFAyJKSWRSzIWtRU/VBTYFB2rnCRyf9D35+7+O79zaX7+W9hAMAAzfDCpjOZodXjsx8Pp8/ePBwtVrnbOboAQ5AjDCSt3VgNuqb3QyJkSgiwg3c0aX6rCB6vZwhHGqBHAFCx04yADQPCKg20OdQ+8UeIwiImj8CBMiIiUiAOUAQqNrvUFAdkVHVQdecbSCq+myPurXupgHhWrz2nJmBO4aDhbqbhzMBMTOnrp103XS5WkUUOAA7vrwHdIcddtjh/7fYEdA77LDDDpcFtFrH4Q1EWvZLYdIxpzyGYSAikQQA4eDuTduIMBGBG2JIkqpPUVVE3Fol1obWiCBhj6BSlImNI0lezfNQhuwYfRAc7nWHe1MGVADcTHJgE2geEcv5goBEuJRcSgEAM6+drRZQTJuUiMiqV0hlzJlFAL0S0E5UM9BZTSu5XLdaOAGE+WjVFxFEEA7mIwEd5tW1Q9VG7e9nzd8DNjmEgFHbO7eSGiAY+38JAUOYhZkImJnHhMcxDL7O2cw9AogowqvEe0PvjbJl33IgW8H3RvocG4a4vj7+uqHpN620o5MGbHZ3tQGpm1cl2O5eueca5VTdwAPJq1xtY7N4aWZa22PzKxiWgNELPCJKKW7OzPPTExKZTmf7h1ewFGGaTCZpMk1Jwjylpu26vF6XnNu2zZaZmZsW2paY1E2IJDWzvb3ZbNavV1oV9iGBRCxE227cr3KHbRnhL0ANfwGW6tchtuLiD79JyWflMc1N1ZwDEWvI2FCGK4eHR0dXwkNVCcmR62Wu7qeLuaqJpFLKw5Pj49OTnLO7LZaLK1eullL6YfAIYVmtltNh6JrOzBbz+d7e4XrdL+bF43MpoJ+J5PzyIgCy+3Epv1iusE1H0akHINW4QAgwM1UELcMwtGmCQm7h4apaci790Pe9IBYRKaVWUuuNTU1LLkUVELNqQRw8TBX6vg9cqc8DF30+zvnBclUCbSSBISDMLc7ufh7hAcjIR/uTt7/28h9897vfefutF5/bb6FvyTqm/cODade2jSBBBKi7arYyROE/+fYbr1w/+Ju//dH/+r//7f9x/zQHDBEltBDqRkUKMRrXbkjcp+8deexN5qu/uJ5Ei18ogiJQZd0FrGM7aLnl9K3XX/jTf/nH/+E///4br97Ki+Ph9MF8MS/DABDEVLIKoSR2Vzerjys1HTRb2Jl6PIAQgyjCSyklZ0kJkdzBVD0ca1xeQD/069V6ve775bKWOYSFED20unCXXACAiYpqfRpiAIRr7jEcIUopOQ/DMNTnfTWTKOrL1aBuAahAIS21ex8dL3/84cN/9w8fLQYDJMSAIKxNNpfncbpFXJAVT2ezwyuHQ86LxbLvB7MID1U7G0PUekJY/SCLwMVTdySA6wivDkjGgjbBOdeKseZNDOEQ5xIqtm94RBN9fp0RgBEESZgEiAOZkAkQwVzd3WsKNIEH0Tgaqvf+cAPAOvwLVQ+zWspQdQgkqm7hJCxJKAk3TZPaBgiDIJSW76333jp5dgdghx122GGHZ4MdAb3DDjvscFnw/f/0X//jf/NffHI1cc7TCTXdLMCDsekaCKRxwmZaFBzCokp2IcDNKQAJhbiKZ6v2mYgiaptyAEJKiZndLFiYiNOE+hIoivLqyy+89PGC//oXvJl7xUYEDAEIqKUw4c3r10nI3Po+DyXnou61URlF6ld75Zd96ybtI4+aUkopSRItWrSM8mBEBHJ3rXy2x6giRgSQqp6qfHrf9zlJHmRYL9wCgh4zvR9z/wzAAxHDghCdAkf7jyqCdq1ewFHqFFd4FC9vFrhhgavyZ6tHfswhizO7UNz+E6NOGyt1AQAQW4oZwqN2JG+F5pstRgBwww0TXidhVVa22YluMfLRflF1dKkmzI/WBx6zeuZe1NzB3VNK3jRh5u5l6FsRRgzVoR+Gvjegfr3eM5eus/CcB3RPKUkrzByqMORSStVBJ0ksiarrKFGtWGBqUOTc5Pkpd9czJInikR+e9C2/QR7zMhUythYcvKnJIKaUWC0gSi4GaG7dZOKqiKRFIwKRPJwCRdIwZABk4aK2Wq2KFmlbACglA0St7CAA15vk6GwTn5N9epTae+Tw4bnFxbY2c4n286/E2vyjfpiBXx3aZc6rYej7Qdq2axIzAwAiNU3LIoDEwkw8nU5ns2mPIUm6SdtNJpKSJBV1QEJmTg01DUdEoDIbwBq5IDnSOnxhdjLkpdmyqAEX9+JhjjVkkBJFgGquvDABvPTC0ddee/Gdb7zxtddffv2lF68edldmvNccJHIGg1BdzDVUCFVzv+6Hfm2qiFhy3l8Nb99oDv74zXdfvvrzj+/90y/u/cNP760jBocCUK0kEJwAicjGrh26mAJ73qnjAvCRC3/zu3/mlf6YGt6vikG88Oa48KIDIiKP3UpuuKl51s4ej0CI5I4RkzY9/9zBd97++nff/eaVabp989obr966mvLig388fXDXhj5UMdzNzc3dEIIR3DSi9mNBAORSPCIIowrhTRMLE9mmmGpqRUstZtdM49SkJjVMVP3Ft11HruruEE5MiJhzVtXqCIEAHiDMCFjyYLZ9WHoAek1fDkRkkTTbk6yazbpuD9tZtLMHH9z74M69rGYQFlDttb6gt9evi6e551ey2IR5MmuvPnd05drR6en8ZLFc9pkktdyoBjAi1SCLTWVbagcYRARwwLZPqyq+t6ONx6D2whFUthoIAaoIvVohRQ2Jze52vvNs/IFwtH7uUtOmBgAsHB0A0CIwwkwx3BghCUCCBAQUEAA88ucBqpaHIaLGbhshirCw1MBtablppGmEEJgwdSl1qVhxxwh/8T/5f+Y/euHXPzY77LDDDjs8W+wI6B122GGHS4RmgD/5q/Vfvo3z5fKoawLIA5gFxgZMCAJCD3cLBXAEAkC0aiFR3QggtLp3ENV5SP3oxiGCmaEaMaeWm2IOGnj71o1bLzyYNeTZt02WG80NAoCpuhkTzWYzZDydLzhLUnOLAELi2kZbOybr1DTCz0RrEWmDUkrOGUb+mSLAPXxs1o4xKfHcnExEPLxt2369XhGVoXf7DDrvjCqOQAxAxyAKJ0R8VL9DRMJ8bgJYnUW25tVwznIDYPP5uMA1jc7PF146J2sOHIknhLEpNbZyo9jMEscvxO0iNr3LWyPNOumv/3qtDFzqxKRfBTPPRQ0IkZrUeKPWr2tLftW9hvt6vS45Azda1N2A6qQ3yD0i2qZlZnCPXDRrnaW6uakRUjOK7AKRUFoiwUeO/uXD5V/Drw5V9UxEMFrNYO0GGIahGYZJSliNfZgR0Syq73BEqKpwapuu53mtDaWUNksbNa3CwkRY5ZnMEUFMLAKIX/EVdfnZ6OJ+EnE/w/1cblXjjPqHTW8HRIwu+RDhDoDVXwkRaCPJ9GrSxOgBxX1wL4iKWADDPQcsAQaPorYym+cyH/LabDC3QPUoHgAUEAEGGACO4JM27c8m1w4P3v3Gy995+7V3vvb67ZtXr+53aCVh31EDpl5y7le5X2kehMJy7vtV7temmSDAHQGOKHU3pzcO2xtHzf6kSZSO+3Lc5+NVv8w6FIcqjt3YcuCZuz+co97wcQQ0nD+8ceFwP+mwP/Em8OS7w6Ps8/nnESJsXBhGY4QgPFvdxDBtm6t7sysH+zeODl6+9dz33v3m77/7jYOWJgKJy+ruvfXJw9OHD2puZ2IZH9imEY4APuYoEBIGQCkaAMAUHtUuQ4gJ0czrs3UYBtVSl1GbpphYRJqUqmHx1uil5GyqAFAv3voBs1If0gAITUPEGCAkyFzDHAICwRlAiAMEkIFTdh/MuNtbKH58svr44fLO8bI4eOAmqu+J+/fLx6/87nq4UJp05erR4dXDbjr5+O7dZd9bQNe2RGLqQDUcub5/1ExXsjjCw2UzCnrywGGbSbGNMjy3cmMxHoIQ3UNVA9EBPsU+148QAAMkIiGOCPPAAHDYXEcxWqNVzXKEh3vAqOaGwIAwK3lABCKieoY00jSJmZlBGm5aaRuhGjjcJmQofQ5wQF7/+J39r//gCx6NHXbYYYcdvjTsCOgddthhh0uElz/Wv3s5BvMyX3Y8zau1ruZtk3jkZbn6Q1RVkfWlZoOf+Q/jpn0xAhBr+nxKiZPA6G5Ro6MYiZAhNY1ZmHuaTV64ceXqIetJlN6rjcUGdV7mw7C+e++uuqZWTk6PzYFIIDAQwoKDgkazZaYaPy4ikliEWUTqlFJEqjkvAFTPie3sJj7d/D7aD7q7u+/txXw+B4jVYmnmtT+zfu6RvRjb+VXU9L+owuLRz/pTk73hjCwe5ctbPfLZapz9/8LrW8IYEQGINl9/tkTCUWW08dWuTtTjdO1cUvxFjvuCgg3H2eMoia5BQHiOzLhkBNZTzePdXd2CmCUZIAAycy55b2+fJQECMENE23btZJJSAnOomWZN0sGHnKUVAESWSAkCtFjGPPQ9izCPvufFA7gFHCr7eG4Nn2afPSrl/lLxa37X5WcyPy9G9/PxbPfI/ZD7vumIhdumIaR+1SNBADBzSgmq3w8AAOzt7T28d2fIAxJduXJl0nX18uHNHUlEAKA6g9eYLCagja/958cTDt9jaK0LL13+w1afKQ/N76j17iiSulaahoUB0MygZtu6WlDOQ7FQVYEILe5ecumpR7ViZh7F3YZh8LIahr7o4E7MmejYbB3QZ12ZroayGopGaIB7FDeHEE4eHq6hCmEc8NyV6dffuP1H3/v2733z9Tdffn6/wWmKlrOWpQ55fqL9aj2s13no89BrHtANzNwNQ8PVrNRINAMsmAKam0ez2d7+m2++/uG945//8t4/vf/LD+8sHpTB6h14ZJ0/1XxzLqsw8NxT6VPqeIynPdBbOvvpz4vHPgS360lROfMwACNEBqDNIxIh9hq8fWP/na+/+e1vfv3rb7xy89rh/rTpGHR18sn9O/d++X6UbHkoQz8Mval1bSvMAJjzEBHEjESAMBp/q6sqELJIFbKau5tVM6va01BKZuGumyBSSm3bdCXnPOQ8ZKLRQ6JJqZlOoUlS/bEwELGbtABQXZtqxbprW5HUJJ9MZ7O9fUfwcDNPBI1w17ZmaEHSToylIA1Bf//TD37wo799/87p6Ro0KhWKT3ZWuSSICEDCtutu3Ly5v78PGOt+rabdpOuaSZIWiQI8cIyArsOLmtpbF7H15zDzx7d0bd4GsKWJz15x92HIANWsmUwt3BXrubU5wTcnb70AGIAc0MZhiwFADbzEaJrUJElMqXa5jDZjrkMxzVYKjoMq7NqmbZvZbNp2bdMkpjqqcuQgRiAgQiEmJotY5qxASbEv+//Vn395h2OHHXbYYYcviB0BvcMOO+xwiYB//uf/23/7n2FQYphOZlT6dek9TAczVQhCIK6WxO6uHghBUUXG4xKImGiccHhgAAa4G0BUa2ZEZGb3GqhHbqbmnrRL/MbLt9c/vXPaL+qn49w0GgFKLg/uP2Dhbtot5nO1AORwrC3Vo2PHOJtDlqoixlF4XDUsSEQ0JlNZICIxb3jhMXAPtwroTXb7+P2IeehLURZhZd14Rm8QT/p5VBoHbiOzLr7hghpoMyn/lFb2PKfwuL9sSOtz64Tbz8DIfcNGCF1DCM/1ZJ/t5W3j7LntvrAdm82B7d7+DC3TpUathQRhGKzXaxj6g66dTKYR3jbN9PCQDg6uHB2t5nMDKCXXfKKiJZcSaqYaHv3Qcx7aJgGAME8mk7ZrSymn88V6vZ5IAiAgfkTIdTn32K/Jdz+TjbpELAwCVt0bhyhiAEwmE5KU2k6Ycy5qSgSqpZQMAMS0Xq1EZDrbY+bjk5O2aWbT2WKxPH543LWT6aTLeVguloioqoTITBHepETMAVBz876srQEY7wfblzbmO7S5MV1mLN3vl/Lxat2WAUppinZNYEOmBcwr54QITZMEqO0mTZM0HImQEBAdobgP4QUAI8iiB16hL92i6BBwfz30EQPgYD4UHcwtwCIc3MAcQF0jDEEnLd+4dvXlWzff+cZr33zz5bdeeeH5q3tXpky6jnW/LqvF8cOyXoPZ0OeSS81IVLOwICLipCUAqJnuEwIhMUsrDUjn0oBMQCavnizfXQ1r9Q8/Of75R3d++v6HH3x895N7D/sCxcPDx0fB5h5+kZg+O8KPO6afusTi3H/P/0rwCC6UJS986rFvs7M3BwQAheG4qkEADcFz1w5u3775tVdfePOlm6/funHtYG/Whi8+OT4uXrKVoaxXphrhKDxt93loTLVNTZJExGrqHghIIoCgqjUUwc2BiJgAwD3MrLZj+fgys1BKklIDCESURLS2WDEjQIAziwgnSRBepfQ19MJUmSmlppQcHrU9orLTSVJKCYjcTVUTQRJuUtNnywrYTgaUVfYf/+z9v/rhT3/4kzv3T9YW4AA+ss/jfy5xRcgDoGma6zeuTybTfj08ePBwPl96QNZiDiwSYRG+Gb/EhfHC5yegN6OhMwLa3QAggmoypKue6Qa2yztX0JcawOyjJgKQUVAIiZBpXGbOBuGhmSCEgsAJgFlSI02SJnGTJDWSGiLyiBKOICTCnIiFWIgBiQi5HcyzY46Y3+onpzuKY4cddtjhMmJ3d95hhx12uFxILkVUpO0mU4oSZem5LzbKX6sSupptVH1vNb6IGAf5CEFMuLF5cDONQIOa3eQ++hKPLsKI5m7m2OK0kbdefen9u6uP7i02dOhmMRAIpEVPT0/3DmYkWErJxdzBrHLeYqOJqleuuWmasVvTRmPGSkAD1F7LULXqB1LfVtUv1UcSNtl9dRNGT0Oiaq/AxEysj9lzj1WBAcCZrePjJl2Pm4Y95n3xyA8XfjvX9fwpjBYbZ3QzgF/Qxp3/6HkB3YUlbn6oTPqW2YjfUvYZ6mngEYgOYeHg6i6H+/urfj1fzOH4eO/atfW6X6/XTsJdUdWkqqWYGQOoqiSZHRx006mbF1U1Cw9CImb3aNu261omCrMaennhWF1SfMWa68uLygLVmEqP6jyjqkWLBlEqhSR1bdsnSY1MJlMiVNX9g4Pj+8Pp6WlIOmobVR2GvmgBBBJxAIsIBPCoxj6INJ1Mc86IPCajfilnx2OOKSIS1poTjs4Il5uCHjyOs76/WByazcwmRdU9kNwczHnTfCPCQKnrWk5imgExCB1RAXJE717qDd+jD1g5zC0sa2/xsM9DhCIW92JePCLAwQPMx4qktS3PJu3tG4ffeOOl77zzte98663Xbt88nAjbyof5sDrJq/mwnM+PH5R+zRFarIYmIjETB5Gktum6vu+ReLa3Xy0AWJI0rbQNkEjTtZO9689lINk7PLz74ORnH/7yb//+x//w3i9+8ouPT5Z6shxOV+t+yEXNNx0qNQovAGD0sR3hjzn0n6pi+sWHS5x7/cJnL54cT+SgN0vflo/H3hwiTMSNSNe2XZtmbXNl0rz2yvNvv/3622+9+srNo6MOh8Xp8uThwwcP+743NQhgwslkEuHM2DWNqppZEkmShFPUCDoPTgkQNo1NYOYASMwB4R5uKikxs6pBABFNJhMRBgwAJEJmCQ+ASCy1iaG2TMWY2RuAISJMtF6vmXnaTVS1Zl2YapgLYB0AIaGbKYAQ8GgKBuph6id5+PB49Zc/fO8vf/izn/7ytEQ4jjV6AITqJIFwWS/DAHAm6bruuWvXUkrz+fz+/Qen87l5qGVCFU2VgIZzAmgYzaMBKwOMVId/TyKgzxfft/WTjSlz2EbEgEiu1Snr8UWWuviNT8q4lJoCjYyE1QXaraYNuoUVxjCiVig10rVNN2naRprEzMiMxAGoHkhIAFLb+yQxUPWAE0htHtSYvXj3oFlfzc9u5++www477PDMsCOgd9hhhx0uFwjooN+LA9OIbnYoPnheWx7cFCGNtr/VBdq0OiFWfwavEuIq5IFRXVI9FuvEjIgYobbKVn2yhzMSJ0aRK/t7r79y+6/+/v0E4ABCBIRWFwoAFI6ulgE8JZlOpzyUks0IPMA3xE0VOTPzVtKHo/kkI43zYiSkkQR31xgj24mqQwLSSFJvYgAjIDwiVIVImJXw3MR8o5P+1ajr81h279GPP0akdkEpffb6p/qsH11IXFQ91lV55M1x4X+fevmiJGu7FpdWM/lULGqtiIQqEUkSMBGmtauZkiRhgWouztUdtDo4Y0qNNQ2U0jStmxOzJMl9hoBawDAzLSU8EJmQmRguOHp/9bvsksuuKy7pSgYAQKiquVVJXi5Dw4yVgWCqYafhFgAeUUpWLWYeAbPZ3vzhgyGrO0hKbdsSQWpSN+mG5VJLyTmnogAgIikJAthYq/j11vcpTv56w6u3lEt7GT+Klep7x6e3Unqpa0zEkItFyUZmXSPmrh45FxQQ0yFjLqWE9+bZ3IJWAWvAApQ9Bi3LXJa5rIsq2uCx0NAwhbBw9XCvd7ogCgonwlnHL714463XX/rD73z9m2++9Nrtm1dmzazSglqCAAAgAElEQVTBFLlfz1fH947vf7JcnA79isLBrZQqvGUSbrtZO5lJarvJbDKdZbVAlKYFQA9wc0nCIrkUNy3LEzQPgJUuW4dXr+/fOPruf/D9b8/X5ZP7x//00/f//Q/+/sfvffzLO6fnTaMCwsEBIi64bXzKbeUpzo0NgxyfpkLPlyfj/A9PWi5CEIQgdElm03baNdeOrrzx2isv33r+lVs3X3v51gs3rl69soe29tXJcHJn8fD+aj5vECf7+0mSRyCSCBHhtpWJEBlJmJmFWGpzjwgDYh6G1CQRWa3WESEpIRMChvu20GLmENF2HYQPuSekCC9F6whGtUiSWr2uo5daxXbXPnoPL6VAxBxPAcDdSylNSkJkuVQuWa24qau5a7gDcA7uQQZM7915+Dfvffh///D9n33ycBmBhIAQ/lQH5RIAAajruoOD/cPDK6WUTz65c+/evcV8rgo18rlQqeMuxPNnCCJRuEMEuG9KEvAky5GzVx+5LeG5bg0iDHdXe8Q57eIa1/IBIAsRAkaYFVdHCDDFcAwnQiEUocTciswmzaRt2ialRIheNHsAYOWbmYUoaMwGgFAzU2+lkSZRM4myRLRIZCv61//9//nr7vIddthhhx2+BOwI6B122GGHy4VWm6FRV7/78ORoNgv1yIpjtykyS0oSNqbLIwJslMKV8lXTXDIRASCgaW09DsBA2iQK1nltwKhOBkBEbYVfuH50tNdOEhQF/7QLRHhUOtoJcTKZEAmTqtUZDqvVgDzdkMlV12wYgECjKSGEe+0PpZp1TiRbqjpi5JKJEICq1oYIYdPESQjolFLSIoWo+sMiACJVreQj+/KLNdM+fmL2BE30Z5Da59moOPfD516xi7TWp2Xdv6VwD1NzVRRIKYEliBj6XkueTGeTyQyIRBIiEXNKSVICprZrPQ9qJimt+vVezhPzehpsqyxuJpLKsC65lJJbt3rqfsZU+TeH3wru4zeJQIqACEcMRGCuRvNAG8mwasl5UDdJMgyDe6TUIDKTiDQijVn4pqBFxElSH2CqGEAIPmr6CMZWDP8SVNBndwkca3Kj0jJiU0f6bbie1f24Hzr3CUIacptyI6kUZTcSBne1GMzGHoRSsnkmCoBwz6YnaqdqA1hvvjbri65V+2IGWCLWZlaNisNHg4BwhECHw73uxrXDN1+5/c03X/nmW6+8cfu5G0fTw1ZtNZ8/XGm/WC1OV4t57telFAuS1LUpJUkiwswI1HRd006YEzFXSai7535NROEx5AEBiKgmLHr4VggbSEDccWpJjvb4RnfwwuT2S/vy0RuvfHx/cf/k9HSxOlmsHp7M56th1ZsDGITDxss/sJZhz6lAawBbfUCMplVQ+5L+P/be5EeyK83y+6Z77zMz9wiPkTOZmUwys3OqQpW6Ww01BGgloPedy/4TBG20VqF3ArSS/gFtJAiQoIU2DW0aaqhKpVaXStmpqq6sSuVYTJLFISJ8MHvv3fsNWtxnHh4kM8kgGcmg0g4B0hnuYf7smdkbzj3f7zzKW7qiK1CDS7ZTwL5eYPmDZW4JgBGEUYRzkvWQv/bKCy89/8yzd29u1sONa5tn79y+df345Hhz/Wg9ZE46tunC60TIw7AmZAjKqeSU1Q0RExNQ3xd9WSAWKHMAuPe1VG8OiAwRrTVtoc3Dq1fpiWZ7eHLur2216m61zhBharXWZf5pWXEk653EZiwEELXO3fw2s/4B7WtF5k57yEMfrdK+BNXaAh0haVS2Sm/cO//Rr97/y1+++7fvnl9MzfZzB9FbNB+yUp7aj2EAxNHR5uTkpJTy4MGD9957f7vdtaYQggD7i6zuqu+XJZABAaK3PXsAgnc/mBDAuyvdq0TdIgCJrv4hfvD0tFy3IGKfTQm3/dL+I851nwmg3pG9vE/QISAcIwh7B2bsp+VkSKnklAiFqFcMIqKHY/T+z/0SCAFCR771ikoCIgAPFqc8Na0QLfjBPRhWT+G5/qCDDjroIICDAX3QQQcd9LTp9/7Zf/av/tv/HFt+r16EAU07Hy8ELAu6Yc5F5Hh/g4p9/BGJgHDpKVQC1YW9HABI+ynW5W6xB5l6rtg99sOYysS3TjY3ruWjFW0vLi2Ay76siAiPznmMkjICIzRWJxZJ2cyatmbN3TuxMcLV4JIT0idqzaFzCANYWHIufarX9qQOd2dmIppnBwARQWJA7IP4YU5I1lqlycwCAqPfk2OAffQs6MfrY3/mN9+UfuR3P5yGjo/688e2ofepUPiye5furuaIrGaIaO4X49jrki7XJFR1t91ysU2E5HQZilfzqq1ZreMu2jHs+TNMstocrUmmcXowj+NuJ2eneXvWplbr3Jc0HlOfKM39afVbeAU/aSb3aVT31PZtZqYKAcfH1zRCVWud3GwoQ8WICFUbhmG1Xoe1CFTV07OzUsq169fu33+wG8e5zgQwjeNut4uIlNJms1mvN7txd3Fxoeqr63ckCTM/md11aQlhz+7F1fDzl8F9BgCPmMzu15CILFIklVRUjcPYLVwsvHqgO7nP7s1tYq6AarFTPWt63trOfVSb1FpENZ/UPMDCq1l01GxEZ1cQeGJapfTKc3e+8/or//4ffPvbX3/5Ky/cEttBvdB724uLs4vzs+3Z2Vxn9xiGlaRVEil5tV6vj4+PRYSIwLwnoSOg1nncXbRWtdWmmpghYhx37o57kJW7d7hwdEIAAAISi0i+du3ardur1++8ZpTPdu2nb7z1t2+/97dvv//TN956652z9x5MNaBFaESEm/tczSACu+WGAIG+B1GB791n6JjjxYOOhZdw+eHtp2wIB4ylSTUCIAiCF7wGEwsT9jfWKvNmyJvN6mhTbp4c/Yf/wT/43nde/8pLz22GXIQozFtr03jx4N6D93daZ4TIwqth2BzfWG+iNRNiYRFTREiEFgZhCF7nSZsSRHhYUzN383DvtiARaNOmiogWZq7CAgCu2p8NLcQSXMxsM21Nm2pr5g4QwikCzL216mYAmLIAwDTNLCw5RTgERsA8z2YGiK21cBeR/no1VW1N28ySSQpImRDe3bY/+3c/+dGvHvzy/bnuoSd+OZv0iPv8RA/4n1FxfHx8cnLCTLvd7t69+7VqOCJiL91dlvkD+lIO9UNNJ5kABIPbQsygRAGB/bVDJCZrERHIHADhBn12AD8IIo+I3uXhqmYWYVd311UPmgA4kLrR727eQWtBCERIHeJMyITroayGYZUzQ2A44XLqR3NmSMLcp12I+hUv0z7kQAxECORAU8DFOI4OAnDtmp+dfQRC/aCDDjrooKdBBwP6oIMOOuipk5op3E+2enB+nuo0nZ7ZeBFtVHdiGfKKiYQ5sZAwcq+WFxHu99sp5R6MYmZJstpsFujzwoAOJDRzMwNAdzcPi+Wi/vk711945sb96UGr5ld8kcs8yfnFRS75xsmt6O324dba3JSZmZgTdwx0v290N1Pr8/KdomBmvQcnIvpE72UisPMTWmud7ufuRJxSaqpNzbthaebuFrqbdh4e1qHIHywW/Lz1KQAFn+Qm9sOP9knufq8mqT/hX3kalVJar1ckkigbs0Zoq6dnZ7dv3yKWOs/gzkylFMolInZn56sTdndVba1G+PWT66UMkTOWIb+TSymqOm53uQxuhoicUslDloxgEF/4Xvrtb8CXw9b8dYoIVfVaOwdazVXbbpqlDOsjFpFaa2s1SRrKEO7nZ+dMbGrjVI/SMAzD39177/TsNCCGoazXazcDhIgoJQ/DCgHneZ7ntl6vUypE6Kaq+pj77bE/gB0rBPvs85fuRRo97pmfeByZl9Y8IgFiQDU3j5kZiTzA3Gf1nUaEt/CLZudNt6qz+axW3RWghauZA/TgMIYjBIQiBAFe35SXn7/7vW+9/r1vvvraK8+drBnrg5/9u1+kqAktk0cAhx+thpNr18qwWh8dEScPjOi0h952a/M0R199dWut1TojoWkbd2MvQ0MIJuo9t4iYS5nr3M9cEQ4RjGgB1X0+ex+ZgTLlVXB59jjdPH75G1/7yv3z6f7FdH87XYzztra5tffvP3jr797/yc/e3M3VI8wgwACQwRgAIPqzRgrY53evgpgu31K9NpBgec+gGSIQQuKgAAZcr/iZO7defuWV68dHiWm33b780gtfeeWlWzdPVqs8JL5zYzNk8Iv3HtybvM2hShAcgRFYW8xVzVr4DpFZEMksEICQiCl6o5/WcGPCaRzbPPX0KRO7e6112u3KMDBTq3Pn1xBR9x1FhAihj15FtFqFRZK0VjsHLNzdrKm2Ws2MeUE/t9YAMec8z9pZJNvtrj1ozJxTTjlpbarad9vSEgEBzCknpg2LcBrSapM3Jz9/9+zBvbd++V5997xVAO0XM/jhz90Tvoj4TFpi8sfXjq5dO9ZqFxfbi4sLRh5KAeT9UMUSkE9JPoDYWALrTEvggICYuPTFDIiIkBQARLQMgeyZKx/Yjk5OM/PlghD5Iy++EIABBVGYBVAQpJcIYwhTEk7MIigEhCCEYdrmCEYhCojocWciJkqJmZc4BaGIiLAQUTiOu3ludVTlYZOPePKoHpBtdXL/v/qff/SEXomDDjrooIM+ow4G9EEHHXTQUyeFKWOJgAhdbY5j3s1tag3NfW7jbjsKcWIppSBh93FFJEnKObEIE3ePYxloFUbq4777W9wIdfVwBHJYGIuOgCR3b19/4dnbf/PG+Q4MHkVF9C92u11O+eT6TWZmlnBtZmoe7s6E0Qc+ARUAws3dHHreKaA3J/bMsi6sVQRYqnGgp2Kbmod5AAAzAGJtzRb4hy8hGuKcs6v1udGPgm88/foybvPnKXc3tQAwVYgoOQ9Hm/tCtVZCSa3CONZaI6K1Ou52xyc2j9O43bXWepulu7ubzbNOdXtxkVJi5v5WMXc1IwQzBaS2H/H+Xd/pH69PR615IkJCSYIiNhkClJxFpOoM0BPQbbPZ1O1prVPTNgxDQNz7uzd3u123rnLO7tZXvHLO0zxDRCnD5mjz9ht/25voVrmUnM2sFELEAKQnlYAGWMKuj6Sen5Z9/ThqEVv392tN04QsUFvGUOEU5hFn7uAuqtVsbjqqmXm12DXdqY1q1b25q7sieIS5B/ZQ6mJAF4brx0d3b5589cW733z15d/79uuvPHf75rXBpvPxXGevwpFZshAzEVIEMItIyim7hbVq5q3VaR4DwMzmceotBX3Cxt2J2d3qPAM4EeUkmJLsm84sEEiQKaJjQICJwM1AESJULRRNOet6dXRcBNP62Vsnk8WuajWvHhbw/oOzX7313l/dvXW+G5v5ri6rqBxACEx8tt1uxx0zqXtVdw/fE3sRMMy1NdNGhCWndSkiMpS8Wa2EqeR04/omEQvitaP87N3br7z88tF6RRi77cXdO7fu3r2zXg1CAK6hYz07vzi/X8ed1hnDKYIAE3G4W1vMXwhgEWLp+esAIBYzq3MDAMBAgDbP2ioCJJGcc3eK66yIjZlq1b5oTbQMq6j24jsUYkRoFh6mDqoNAEQS9go5wYTEEcKd9Q+iioipFA9HwJTLuBunaco5l5JTzqbq5gGBRNzz3wSIkESEE0nmPLgMM+R3fvr+j3757ltn03n17j4/uhb5lMA3Pjyq8shKc+eVbTab9XqtrU3jVOeaJBGlK4SWxbmN8L0BjVcfy5yjX0hhMHNK0mEal9WC+8P/MmX1QQAHIhGpakTdT2382vMFIwqxkDCAIGVhiiAIZkpEiUkIhVEQEYI8IiyAerB/ySR0ohYKAoaDQ2i4m7Z9i3PT1twa4GYtAOiIFnbz2386vfPip38dDjrooIMOesI6GNAHHXTQQU+d/uN/9l/+b//9P5fw6xt54e4z4zrPZ5t5e7ar08V2d3Z67u5qltSbtqq1z0WKLO09qtr7CIlIUko5Y0LihaV7We8THrjwVcMiAhN43Ll17YXn7ib5JSEy7hmPV/DD4zgl2QFAzhmQdz6qOSLWWt3d0XsWhwh6/yHvvcJeu3U5SjnPc7d7WmtXqtWxB7Qv4zzYEY0A/X87BjDch1K0NuuDo1/AS/S4+sDt5a/b5E/hfH3hwd6P1MeTH0xtnucwA0SPQAhJXEp2cwRgFg/Y7cbO4+g2orZmZoSISWIXiEiSiAhmVTVtGtn7goaZt9bI3dR6vPCT+QufIur+/wPFh4yPp+LpXzJt902mYGY555QLEampqi3LYBGqSizMxEwB6OG77Q6RmMXMpmlqquFWW1VVVZunqR8nPVxEmKn7kx1F//ibCZ9wp3UP+nEe/6lTADT3d3ajBwQgaSuMM5FIeMR5VfAgwLnZrG1uzSKqxdS6OevqoRAK+87ciNhTGQCCMI6LvP7S3X/4B9/7+7//rde/+sLdk/W8Ox0v7tm0OxrS3ZMX1iVnYQb0iD4SMY3jtBt3F7tptx23FwCurU7Tri8nVK2ETMQeSMwioqYewUR9sVMDhJhSzpxVfW6ah01i1mYQwESDCIKFtVKym+12WwuAcKijmZHMq/XxOqcbRVZHx2W9Keu1Bpxvp1++9Xdnu3FX2/v3z3fj1Jp2Hkgp5ee/+MWv3nqTJI2tbcepmVtEAJEkAvKmF6en4/Y8C59cP75z+9bJ8eburZsvPvfcakgn14+/8sorm1XJgtc2m81qWA3FWtU2m9bd9nx78eDirfM2TzaP0+6i1clNvSlCDDmZaqutU3oZYRonV2Mi7sNHIg5oDgZQ1efZVusjlqSqGEEhEYZBBIxEnFPm0k/ZuazVTN0vJ6aaaacqIYuIFBlUtaoiZxFJpYB5p29LbwKVJQHt7gGAhAAoIkdHx/M8T9O8Wq36mFevOwZAEWLGCOVOdUAKIHPCPJxN9tO37/8/P3nzT37w44uIiuAfHFd4Sj6JVzfj8rD3yIGFiEpJ69Wq5FxbbXN1i5xyQMek9yroYE79CjA8CFFEELAXb0QEef/EuLr2DDsSBoWHExEh7htBsFvYHzhSEVFKCQC16Z4V80FdssqFOREnYoFOdhaKQHcExwgw7xd0LNQrqTuXyM0QqC9aEDEhRVA4BIJpmDW15ro8CRJKJQ/Xrh8dnzgBVUXA8x9/7/i1H37eL9BBBx100EGfmw4G9EEHHXTQ06iZr2OeZq0XUxVOOWf0IQiJZT2shZg77M/dTGtPMAFc+svLXR8iMRMTCkpKqeScc0qJe954aadBJCIRoASch+Mb713ojWv5bJ5qe3iD8dDAQ+ih1FyGYSitqUcguQgHgD9kdQSzM9ueIr3Qe23pGgKR1LGRiPxoQdxSs0Q9CAYQsXx3+UYAIokIC5NyhH15/JzPcUOfTt+56xNtm0eYOQQwswe21sJqSsmadWcZJLXWEkMfwTVVREIEIkaAiBAWzolzZkeWNI3jOmciRCQIcHckBHdQoysNXb/mNbi6zfFRf/ikdZUS/nn93k9tJT8VHnRnh4YZEzYIbS2zlNUgKTELIE3zFADEDEC1NuRIKedcalM3H8cJiVh4nubddtdxQeM4bi+2OeVOpXf3Os8d+Lv8Tn/cJ/7F76jfviJidj9rLe1GditMlYjVPOC8VmhETWvTatasI56jqnU4sgZ4B1uARwQGEHRobDx/5+TVl+5+95tf//bXv/KNV1955sbx8VrYdikaJnIe3KzOtdWK0U9D2mqd56mOU5sruoIrmA5DFmYEZCTuEhZJxAJAAZDzwCJAGO4BQUwiiVnm2gBQJAWgA3SLnAGHJBjursIIEcNQVA0Ah2GY5jq3uhZjRnXA8VTbNnYliFLAC9fys9dXBrS9e0MtiBgiIFzdv/ny7Wn+Th5WwGIATU09HDFJRiCd67i9mHc7RlivyvHR0SrJkGXIKTEm4cyNtaHGxfbeRTiCh7m2edrtwtVUp2nnphiGbhncMRRC1cbaksgqFTODMAhfDwMBEkSvAcwlI7EBzmrMLhxAQITHx8cYju4A3q8aSs4IaG7dLZQkPUVrbg/TshBEXEpJKRFhrXWeKxEyUz+wL/1yy2WI9IsEiKi1bXc7Fu5/cRhKSol5AWh3q1rVa60RBqiwkD4IgA3Szsf/91fv/cs//fN/++NfXAQ05IC4whL7UujhsWUYyp07t65dOwq3X73xxttvv316/wFJBuRwcLAIBwhEBuz9zNCdfQDouDOAcLfobQkU/YOxTAWoIjMChntHZeyX4h4VLh2/2tS09Z/5wLZ245wACJCQEJECwEPnRuEITgjEBMDIhIHhYO4IgUyAEQhBS7t0Dx/Mtan2qIEjAhMJS8qJOOchl9WQN0fDkLdtNkIktt21P/qjJ//KHHTQQQcd9Gl1MKAPOuigg55GNRruzc+9An91frG7tSlsA4YCU7YCgb06qbXW/eBpnns4lJn7/duSgO6pY0KPAPcwB3f0SIl6EhmXnAlzSiQJObXgZ++c3Lm5efd83NYKAIEfxOd6+DhN683RUNI8i4ejOQIGYCyoj2XUmYhgaT6ECOgEZ7hs4kICJEJyd+t8aghcem9iT+foY8mLf93jzn1Gs/sKZtophr/d1+egzyoRGVYrTMnMiQkRx3EK86bq86zaQDjnDK5E5O737t27duNmX3EBNWYGAKuzzjMGJZFOt+yp+ZRSTomYBSlq9dr8EaT5b9AX4j4/OX3ASv5wMv0p/eDsWUELA6GPU6xWq9q06Y6IN0fXVsPq3um93W4rw/FqtbaIWus8NyQehvXJyY06b1ttTdtRuQ4AwiIpAYC2dnR0lHPuv+L09PTkhIWlFOwRvy/ymX8ZFAAasWsKMaWIQbgSMZtHjLUFAjbqaCbzcAAPMDcFsF6lB73bzxGCEYrQZsg3rx9/57WX/uDbr/7+t77xlReeuXX9CKxa287zVtvspoCgTWttaguxotbaWp8Caq4qGIkolaGsVggBSDkXFo4IFuEkROQO7l7KSiQhgblBOAtHgJknQmIuJauauQeTm2NEYgRHcyAAJGRKQoQAicnQNRrpiM5k3sw9AImRmUSGMpAUJNkMgUiSEgK429zqs5tj4ht5WEkuJNLULMABO4bCqrY6a60YzkRJmAHA1VoliPB5OntQwwN8Gnd1nlUrAbraNO6YkBDVGgIwoQgDBLgjIhOpOyKxCBIBJEIQIkZiiH45kLIAcSANyyUDVAtiWa82i2WI4O4QMZSCgKoNEJlYkrAwES4jTUSttV4tmHISEUDMKZWUiHtlMogwEUb4kv8GQwimfqI304oQhlCn6KtETd3M3NxyRiJtptbMNdAi3MPDEbhgWv/snfM//9HP//j/+stf3J9rYBAH+qNFxR8+9D09H/wPbEkMQ7n7zO3NZqXW3nnnnQf3H8zzxA6I7AERFuDQ6c69V+PRv09LrtwwAhAhsC8Ad6wZhIcaAGI4EAFSuPelfoCHUI7eoeruYbb/gQ+mpAOAAIUwEQsSdgRLhJsDBGMQIQYiIAEiUCecR4Q7EGEguEf/KLgZAnq4aXVTZspZck4lp5xEEpXVUDbrYb2JknTeAQCm2Wt5gi/LQQcddNBBn1kHA/qggw466GnUud24Az83iLFWun6NywpDxfNSrKTNXB2cSZhkIPScTK0zGVubVdXNiVBEOLhpm9x6biiJlFxyTilJjyABIgBxEimDGg9CLzxz+617473zat0kuNpzHqBmF+cXx8fHx9ePS+EAIfUel1n61sFVQyMCgNPiiffbFRFGRCI0i31mBwNctS5Dt/So10wP25jczd0IkfsWEzEzkkC/c/8CrLQvgZH3xeljbuYRgBAZoM7VpwnMUpJRteRCpSBATPNut0U3KXG0Pn7xxRe5DPrOOzqOCMHMF7ttMAZySkPPO6eUAGC73TbVuVZm1nDIJeDC3fwT0Vq+KA/i8zW+r45vf/gBP3Y3PB1vZkRmopRsMkTIJXvEOI0kaR1Lpl2EV+tVKaWpzq2ySC6pNZ+nOYkkSf1dcfPmzWEYTJswl1JazuM4nXiICBIdHR+vVitmjlAze8wn/7t7EKhu2jwhzRB1WkwudQskoOiEftuvSVqvQQMM5ACDCAoQhEJw64i/9uLNf/SHv/f3v/P6t159YSWEvt2+e28cd7XO4TrXudXmAMyJWXp/ACJ5AEseVhuIgAgmyCIlS8mJAI6brldFmOd5RiIiam02M1gOBBFmbZ7cfbUe5mnc7XaJEzNP89Y9AiAQWm3hjquNq9V5KqUQopplEUTYnp46OALuzu4DLO157hHYkQboi6Hm3reYqK8I9Y4G6CdfJEDaH536+ivQHjsDHmZmquEO7hFOuIwFdUiumTVtrbWUEhGhh2kYABLuU66k2nZTG8pQ1nlFZGbVXXIZhmEYhjZXcE8sR0dHQxnM1CMCMZfCwoDYmV6ddyFM3VH0MCF2s3mcYL/GzIxE6ISmZq1Gq+4B1GzGgFB1RGAm7Y/glktCjGkaa621VVOTJKWU1po2bWoAQEiMjOF9BVvVtFlncCBSIHi4hgV20xq4bOSI/vwv/uZP/+Jnb95vY0NECiTwjnm5qqtr63g5p/XkPzq/WYRLayNcrsSVId+5czMXaW26uDhTaylnSQmRAxDAo0+KBcRCLNr/AxAQTBgRqsZMTAR9+qD71QiIqE09Iol4uLsHE8DV00iHMyMzmpl2+zmufBeXbcUAJiwkJaUEBM0AEAEZUIgSESdkJEZEWIoG+yO4GwYEYLPmTd2auxFCLiknKatytFmv18N6yMLAhERQhlLWJV87uj/prlUA1vHkJ+/+8rf5Uh100EEHHfS4OhjQBx100EFPo77//e//7//jPzcAdeJcGFZad4gkxMwWwj1kDIHhEBCEmCSJSEDUumqtmRougVBKqubWe9jAoo5TmydEuBzV7HOXwGTpyOp06+RosxrwI0G+CGZ6dnZ64+YJAnj02U/YYxuDaVFKSSREBPbwjUsyNQBaLyFEQCAPzynB3lPu8A2P5Zb8khUK3Srv+WrzMgy827W23N1/0XoqqK3Bcr4AACAASURBVAVfJiFgeNRZhEczr61EzNMc1ApJAGBKkjJo61DelDIx98w+htc2r483pZSUM6Xc3ypNtbYWxJISS2ImIgZz0+b+CRPQj6XPK0P35N48v5235eeIDfmg+hyEu2ttrTZJPKyGnLOpXWzP3U1YiMhUEwsjIgAisNB23O7GXZiB+/bi4s7tZ4AEiQNgnKbbIgHQWlNTbW2apmmem9qHxs4P+rUKAIsA8DBwUAIEBAsHCPBw2PedAfQGwFgA28t/M8ed60dfef6Zb7/24t979cXXX3n+uRubbHObRq1za80XaGwMKZWUkJg5sSREJCYhadb6qipEQEDvwAUI6CdHoHlqU0zaGiwM8Rbu4OEdARKuWs21zVs1VVVKbg1UlYiWnC8gAm3Pz/qjmmr3hSf3JQQKCBDmBgBEpE3dHTqlGECtLfz5vgF91zykWS0+Y0fvBoBbLL7zwqag5fea98zww/VYAGJmEGJglMwokpIkIfalghhJuOeO1ayUknJKKYkkM+3zUiWXXIaZONwTMYkYxFSbufWPSaeXmHkfQQAEJIhlqgkRwtTqPHeDEhdb2bEvIHf0MGB49MknkdQzsyyCCAE+z+zh8zz2J1VrNdM+KeUebg4BHqruPXI+jaOqOQBz76Bkj2imu3nGJHlY5/Xm3kX92U9/9MMfv/Gztx6cN29B0MuaA+ODx8MPl/59gcIr6OfeF93HxSDncv3a8TPP3EXE3W5nbjlnosRSkHjvU/eP4sOzXCz/6p+JpYVzqfcDiB6YXmLv1OMLxNSH6vrF5SU9DWOZbLPW3Kw/4MNmhUcx+P0lR/N+iu8F0/ucA/RyQUTyCO3XbhFupm1mDBYkBmFMSZhSzrJaDSVLKXmzGYYhlcQEwQTClEtKJQFC0+phDvRf/4t/8Q++/vXfyot10EEHHXTQp9TBgD7ooIMOekq1g2vHtFuwt3kNdAoRFI6IIIIYAGDqphbhEcFIpRQkLCVra6rqqu4R4cyLYW2q2lRV29z6XWi/dUdGh6huslYwuXvz+vWjlTBYn5d+9NbMzC+2F7txN9e5zrVVtSCznpoCRKHgTkhAxF4Z1Itx+mRu5xKq7ovXAwDAA4hQmCUlZiYkj+WfPnIbEcTdewxV1Vq7fb292Lob+BeSgD7oN+jjTMkIcAfTMvAMsEzdursvkG8QZuZwRxZmCehwcwv3MNdaATa5lJSzuqk170BThJQTEDkgERMhWOuT3YhxxX64XF35yGWWT/gEH/9Zf4Q+Dk/92PrCnZTPQT2L6LY4IWauTSOCuTPA3V17RtDNzIyICdGbgocII6G6mlZGAOY6V2saEHsiEHbrys3UbDEj/ZIDcDiSPIYsIsDdghBhT2ECCAePwEu7tTMAAoAQRGhIw51rw2svP/+H3/3mv/fdb7z2ynNHGXw8r7vTNo/uCgA5ZaIc4SyJRYh7By3llJiZiZo2NevzMt2A1tbm2kxbmJHDWCdttYc9l1f20jhbHDkzb7VO/VSlqGY2T5NIb1MwkUyE81wRgJnMDACJeR4nNxuGAoDurloRkYV7yQHv/fZW67KqCggAHt4NZ4Cevl1o9eHOxAEB7owMiOYOgRSMhEiYSDow+cqOD2JhEdgX9jJLYkkp9fMmIBAzMUOEueuQAXvdXzJnN0MAYUoEzmQRAFHr7O7b7VbNwl3VEDElhgDrBZ5m5h4eSMjE/eMZ4eGGEESsqmoq1BPg1EspmqqpAuJ6tQIAcxcWIkQCn0JNW6spZRH2AGvamkpK4dGaAgC4W2s5JSauTc0DRYgYWIjIzR3QAoULDUdejt5+880/+cFf/+iN83fOpgnAF0f36nH+1339BQqvGtCXHyIAQMTNZn3jxo1bt2+9//77p6dnqtYrG4lzB25c/rDDUtq8D/kvh7I+gkZE3axeMGf7fUJEkXpGH/ZXa+Z7HD4CIHh/kMl0+YuXn6Mr7vP+CQQCgDshCCAjEAJBH58Lj+g59DAFCARyNzPzNjNBMi6DSMmbzVCyrIay2QwpcU5cVikJCQMDCqEw5SwoNLvWaQwHZ/in//h7/8MfHxoIDzrooIOeah0M6IMOOuigp1QGwy/0+a/LL7bzfHK8HtbX5t1FU8MeMdvbwsS03mzCvTU93160puFuppdes7kRYb93Z2ZJkko2bWbGHQMNYOHNTFRpGGIoX3sl//gXb/74p/DeDia7BAACQL83cgA4Ozt/++23W9WlqKkPfiKHA3NIYiJeiIER+1Q0wf7n+jiyiCygUAgEJCYmBHeLDvXA3lIUSIhopq6GvWaOCBBTTmUoZmqmB9foKdPH3dLvI3IULoiOiI45ZwvIpeScQ03VICKTSCqA6N0kdCcPDJjnGRAJUedRXYEQmTklTqmpNXdaBoMbYTxMRz66EVe+eCwP4je82z6jo/EE08QfzKo98kvhU/3eJ/ipiwjvY+URAIDEIlKt1VpTrrlIyVlHmq2aOaGEW5saWiBhM5WcRCgxCdKQsjbtLjMiDKthQR8QB6IIlyGnJIgan+YZ/a4ferxP8y9vHwSIQO+hTFxMNCBCd0DwjPDcreuvvvzCP/z97373m69+/ZXnC7mgtqrCPByfbK6dcGdLMYV7naYAD3dttc7bVuucJNzbPBFRBPSmOwhADG1NW0vCjEiAdZpUGzH3EG7fGozlJAQBZqqmEYjMANw0zMAhWQgiOYoZoDvnQdWmaRZmRFQNSoUTRp/JgEDkPmJEJMzELIutXDItbXsEABTBwkyXPnLPZZua4f7s3FEeDtF7DkREJAmLPcIQCsDe8dCLFIiZ+94mQHcztwBnRKJorYU1UlUzda8A/erATHPO6/Vmnmutda6NmABinmtrzTRWwwqJpnPPJRORN221qXvJBR20NXVjltVqg93YdN+I9CVn6Q0Nqu6dxdJXAFxERGSeezkltHlWC8A8zzZOjZjNVJuuBjT37Xa3PGE3wpmIkiQaMuYSzEEIhAQx0Pp42NDquEL+4Y9/+a//+s1/+/MHDyar+xRwhGO/ZML4EGGD4GlUXIbrifD27Vt37txeDavTB6dvvvnW2em5OzJnIAUgCIyH0We8vMK6bCBc1nWX4TOACNrDRmKfgF4aFACICQG1Y1hg/4jgAODuZuZuC+rj6nFv7z4TQCJeSy4oGbkIcd/5CA5hYVArROCyLhARQQDMVFZ5VfKm5FJktcqbVS4lpcRJUARFgkExABxLWQlzLy+11nbzZFqL0Fzlq8+d/HZfpoMOOuiggx5bBwP6oIMOOugp1anffAbfbArv3nsAALm2eaqhM2MQARHC3otl5ggCRHPrQ7vQw32qrTVV7bRliABEB6DOo2Ti3hnElADZHVuDlInLs3nzwrM3nr19fPHWbu4Tlw/Vb/ahznXcjZvNkXlsd6NIIhImAQRzt9lo2bAgItlHw2B/e6S9Ry6iznXpLEKEK73t7t5Bz95zNojm6u6E6P27iO5eSpmn6bf+4hz064RX/v2bFBEW7gTjuMPwxJmj5TxMTZkSA0FtrSl3FwuJkIMcAYacymo9jqMbmEVPWOZcUi5AbA7kUbWt1kcpSUR40+i56Y9BcDxR5/exfu9n2ZIvPMr3uQn309o9ncolM9M8zoWZWAjx/OwcIzZHx7kM5+cXqzIQSWvaWl2t1wCAgT34PJSSc1ZTAHBzMyurYbVZgeSSi5t1dKkwE3E89j484Hd6thHg6r5YKMqB0IvI4No63by++epLz33z1a985/WvvfbKC8/fuXFtnUNnr+rNI1zDHUHNKji4m9Y6jQiB4GGmrZq2NoWr1nlike5BR3jHC9Rap2lMIoLUa9cAEDtTF8HMHAKBkGhffSCJ2d05pZREzTnBgEwsAaimRCQszOzmqkp7d68fTFJKgBARC2EeIQKIiEVo/2OXZ72+b4QZ6RHTs/uD/Wd6YBkuvdJYssbEEtR7eqHvZYQI09YUARgpxLVVd+v7yUwjHBEYqV8DaFMECAhVWzKs7t6azrN5mFkzJWIiYkLOGRKJJCKGhCKCiElktVoDkjDHsuoQSMgiy0pfRE9775/snrxAbNrMtDvjHbERAAHkAH2H9SecS0EA9yAiiSDOPWpLABGGAMOw5jJAyh6OAIJBIlyG4fjm2w92f/3Lt/+Pv/zZD3/69jvb1gLsIYZi6ah4ivXhA8ji8DLTrVs3r12/Pk319PT89PS8NTMLRCeRbkA7xp5y09dY8JIDHZ0Xvk9E79++cNmzsTegHSKICRUDoKMx9gfCjteGPkJn5hC+hBLwYfga9uceJk6SyGEZiIjoZZYRC8Qc3BEi98ZKoiSckwwlb0rZlJwTr4oMQ8qZRRDRhSERCEWHgfSIuDZFRwWoVcPAAY9vwbx7OpcTDjrooIMOeqiDAX3QQQcd9JTq+9///r/6n/4L0/H+hWurJ9xs2rJrJpDEmJiWPj/qN/4icnR8vARgAAAgzFtrtc61VrVmZq227kl3XIaCAYIgS8oYEMROwiJ5s3r+7o0Xn7v9xvtvnU3Wr/i7Lk08N3O1k+vXm9rF+ZYzdWyfuavWaRoRqZfCMXNEmue5tQbdD0A0U2ZOKc3jZGq4j8/1GA4gXnUM+9AyYnc3Aq84RDlnYt7Prv6u20BftD6p+wzL3WwD12mexQMQ1V1EbJpbrxSUlMow7y7EjZiB2dXmqeo4RTJzN0ckTqu1Es9Nt9O0Wq17a6UFbKdxQ2tmAQDGZVXj4zbqc/SgH+uhPi8P+rPErj/FIzzZjxsiijARAzKQBNDcnLgEcVULsGF9dHF6b96O+QhObt4Yt7vmZoDAmdOAlAPEgltrD87Pj2/M7r6bprPtxThP59uL1TRisnHcuWqbxjpOOlu446d5XoeDzyU3gPb/0wPHwYhMwITP3Tr+9msv/Uf/+B/94fe+9Y2vvmzTRd2dzefvliSZoILO8zzPk7m2Otc6W52tVWuzMApzlt4PENqqW3OzMGaWlHN32IgwwppWN60BYZ5TzjkzCxB5gHZaMQkgAVHnSxCRmqWcUs6tKRMPqxUSu8c0TcMwlFJC+3oqtdoQIKU0TXOED6tVB+YSETEjYZ2bB4hIGUqf71HVntFGwH3l76LlTdOdQITuccfeiW7aaq1qpuoIrTctPAylBrR5mucR3AhRWOZ5VG3goNZMm4f3isNuAJpaKYWIWm0sLEmYRJvuthechJlFUo9cl5JzHkTSPFciXg2DmUc4Ig3rVc6ldv4VMxGq2W4cfQ+LMHc3D3dV1dYu57TGcax1wqWCEUopLAn7zAoRdWo/0zCs+us1TRMgDENxN4Bgos6GzmXAVIJTrc1dGTyvNrw6xtX1X/747X/5r3/wf/7F375970LxYSvxfvAlrhCWn07Fh74ORBDhm7durdfr+/cfnJ2dj+MU0VPzmgOQOAADvL8EC9v8EjgDAFeWTPYlhNxX+Jd3UzegzRBBIvlS5nFl7G0/xxDunQG9X2tCJIqwDxz5kJCYwszcDD1czVVNAZx64BqAEFhoGPJQcsmpJMkiq5xWOWXGnCgnSgxEgRhCKASyh4y4WajVafYkwamZOzJi1PNWjtOTfIEOOuiggw76HHQwoA866KCDnl4Zwfbo5vDue62OsMlmbd6e7dqO+o04UhnWuaxJUo8Mb9YbYXY3ZmZiEk6EJJxK6jcbqqbatNbeO98JzGbmUdVjaq35DDwNm7h5NLz07O0f/M17DBMA2j7gdqlpmk9Pz25e7NR8HHe1zsSJOfXUi1lz990ullJBxNaamXd/sG9tSqmUUrvfuA98dRDhlezY/l4IoONCzOzSnMMFNUkpZ22t5+CubOPvuiX029VjuM8IkIRLyQhBSERsDrVqBNVmR0CScmCHOLNa1FnBe7xOWkBrhsSwt2/Ao9amaiJJUlYLANRm81xr7fWDsM+Afb5PFj6/99hHJuB+3S/9SH3YA/3kbstnfzqfETzyUULADi1dMAXOLBhGyAAYiJJTLsM4Tq1pALBwygWILAKR1aKpq0UgccoOEIQp5/VmA7EUl1Kv8PLIKaeUASZt+vi74HCcuRReYZgs8efrm/LC3Zt/77WXf++br377tZdfuHtjTdO7P/2LqKO32XW+MDVt81xdNcIIofcVpCQloZMgACFQBJg6uGAYQoS1uTUi9wAk82hTVQuUdVmtELDNM6VMuXDOyIzI+QiRmWQpvBXmAI1wWhr/sJORiTjCKXwjAwK6VUJ0U6uOgEgU3oTBPKZx22o1W7xdiKi19lkfEemrX2bWz1l7HsSCpOaF5tF6OwIuMfElTI3M5u5mHUWFiBHgHvtBomCgCI+wiGAiZkYi5hIUhIxUUk4AaPtBou7z9tPxZXw7IlQbEXfAUQQAEDMBsSFRoojYzg06vyi8nl9EnM/dgEastfa1QofwvRGPRNpafyAMTyLDUJiPIlaSuMNYeqNsIJla/0lhJqQe1Z7q6BCEZI5ZmBDNWqJAgvCKGgRREFrEPE1SjrYX87/5s3/zx//3X//gr3714KIzw3D/TsS4umD9FLQVf0IhQgSsVuXmrRvXrx8j4bvvvP/++w/OTi8CMIAAqekV5jNGIDAyIgH0Nsj9FMKyOh+9s9rCw/doo/C+3NF/0swAsSf5Yz+UBhAdwRHu3uEb+6LMiIcf936txkgQUc0E3MObOYZBGEIkhESckySRLDwUGbKUnLKQMAlG4cgcTIDgEYHQmeYZISBMm3fXfNxOfSvKkMu1Qb0hQExMef6j/+ZPvpAX66CDDjrooE+ugwF90EEHHfT0asqrcnaaKAAjlcRtNdetqRM4BLhjq+SBgLVP0Zo5E2mrna4hItRDV7TEoiUxC5ece7XRQwGBGbsFBhAw2M1r6xefvX19k9+7j5OBxwIXvPTxVHWa5mmaRWS1GiKASFhy9yCEWa2p6hWQpSwVc706zD3nvFqtiKqqujkQ4sLnBAR0XziDC65zf+tIeyRIxELJHHwAADML+yQu3kFPTp/UfwwAIkrMYJYIEVEBPDostPsRAgFELFIASNUWagxxBGh/H3WGL2CoRYCZE3GSrF57h5iqNVMkDFzutp/ok3/y+hwD2l+GxO7Szxbu0dS0NkDUppJy98uaan9TRHirlZkBAQgZkYlMO1oeIYiIkZgRUy65rKy2PbCUIgCQS1kLZ4/J3D/bRj/NEcsnLXz0Kzw62jxz6+bLz978+kt3vvvq86+9/NyLd68nqPX09PT0XmhFV4IOizLr5i8iMiEERXAgISPBApUKW6rPuJ9EkJmBBIlZEiNBUwYklmE1MHGYMwsz80KEZmJGYiDuA0BEqIbhLRA0PJpDZ0W7QzghsrCrhTkTWdP+HhMRFrbuHDdTbe5uWgnR3VutqubuIr2Jd2nf7ZZdR/G6u4f3Cab+3FWNiJCQENUsPJB5QYv0CGsnjXiYdbucmAXCI2zfTLgs1wUAkANASjk6D6vzuYmBKIhApPd2RiAAOiXrnAtHIgYgrQaohB3z4e62hNk9+om41tad3NoqwFL6SgiBwMwiTP3wnnO4CdFQSv8gpsQ97y0igWDuKBgBxMCCCGG1TvM4T5OIMDOEhhFBmCoB9EM6ICNnB24W41Tf277zxv3xf/2zH/3wJ2/+6r2zFuCIgAxLVcY+AI1fhiPeorhMya/X67t3bx0drd39/Xv357kSCUliFiTZk0wAIGAxoIWQIsAtfJ9xXuziiNiv4vserB+una4fEZccG0B8pMKwL5lcetbQ3fH9xu73a78+ZEQEcO9UNQgCChTgRFSICmHueefEWahkHpIkQSEkiETACELABAsix90Nws1d3fuFX6gaBDCzBWhERWwBw/reD39+QLEddNBBB30JdDCgDzrooIOeXv2Tf/Kf/C//3X9KfLJmXg+rPGQrYWPqNwgGMFUfZ6utqZm773ZbU21z7eTllFNKKee0Gob/j713aZLkurP8/q973T0f9UABVQABNNmcZk/3TLdJizG9bEzW+hI0m0+gryCTZLJeaCPZbGaltRaakdmYTAtppdFr0a3uoTVJiewmATZJAASKqEdW5TMi3O/9P7S4HlFZKBAAgSqgCvRjMENmVqZ7RLhHuN9zz/0dYnTzlFPX9cMwDBAijNslsEhY1dI4AVIgBeBL1w7eePXlV652d+5jWXmzBojIHidjqOr+/v4bb7xuFkjS9Xu1WK0VwGstpU4A0Pf91atXAUDVNptN44a4e+76vf2Di4uL9Xo9jWPKOYm0FcoRYWaNjJmyIIKqxqP8TRuLanuaYzcS0Wa9vrTSdtHzrobg8FIg3NTMHZDHqoEURAYBAQYYwIAcSN6iVQrFgCPWU000gHRB2XwNlMZJq3o0p0myB0GAI2KWCqDRMq9PMbkcj3/x5Zx1lx/2k9SO30pPPcT9lBURpu7mVb0F9aZapnHinMzNAcdx0mmMQCJulaqbafSIlHuanWUCZHMrkxIKE7nGZj2VSQ8OUwSpebFwSo5p0hiLWdBvn5Kcc4LLJ0/TDgP1jVu3/ul/+O/96Xe++c2bh/twwdP53V/e8bIGm8CLlYphwsiSRFKfpOV0k3CAqzkEqKqHAyAEtssBIZo7AAbKcLCfUucBfT/kbmjzDY1cm1M+2NuPCHObq3g9iMg8apnauh/V4l49qmrVWl0NIdy11pJEckoppbAIdyGqpYybsWGjupxX69U0lXYBZWatBQDCYyqTmyFRlzMzq2qpVVVFBAIahbx50OEBEMwSAOHhQRQUiC31zDRnTGFe52EQs+/c567rctf10zSN46ZFrYlkvvghsbTuTmgc32paJ3V3mZHZ0TzxtjQEAdQMIohwb9gXTuvNGiBEmJiZWYRUi5lhRN/3OeUMGO4AkPvcktU555SkccBaspuIRKSW4qbzSiYEZmpAMDc313Ea53lBRESCgDKN0ziWUoZhaODpMo1uykgtA16rmkEAGYpRMso//OlbP3j7/R99cP5w1BJg0Kz4FFYhLk0mvTDZ59lSbl7/wcH+a6+9Ogz9+cXq5OSERa69dKPr94gEAKZaPBwa8AZb3hsBMHy3nmw2oGPLiG43ewDeENGmCgCSkqm1APu2rhDdZwvbzEyL1rq1gD9eiEDYZiIQIhAJhQQlAWSi/ZQzQSIQxiSYGBmDERJhJkqMjMiMhMEsIiSJEKLUWlYThEE4gDe6ek65TQJR7szRgBzgz//1T/7sH73yJRyeRYsWLVr0BbUY0IsWLVr0XKtSOaW/24s/Pjo9vXlwwJIwZSIABAciDsngQS3hsxnXtZbwMHdoxgxTCwa6e4DXWsx0HNda53hyGysiYiAEIKckQsxyVfqbN+L3Xrv566P18eqkreC02QKYO9fdbLVaHRzs37jy0unpWa0FKbVSIXMXEUkcETnnndNtNsM03V1SIgRh6ruUWh8NzbVjcAl3SYQAYdIiNYCILRrpbjOvA7BMhUXcWt0itJKm59VY+1pqh9fcmXGf/icWOBY7N9ucj+P5xko5PV4BYj/B+RTZ4eGqrM8uuBv8IC4mRIKN8do4VB+clz0eVlPsKY6RHl6Uhyt9sNKrKx2L3TnZ3DkdJVG3qgejXUxetE1ePMVzAj/Nev5YIMZnf30+VZ/seH72N8Bz+lZBopQSBJr63v6h7B2er87T3l5xXG1qv5f3r107f+gXFyuZqgLppMC5Bo2bQpMeUjpbTacXk4gADyjdVOvFppyer1dn56/93h/0w+GE6JxXCndPz/rI52NZj+OLn5R/DhQBGOvVxa9v/+o7r19Hy6FrmFZY12QFIZCZU6uXAyAJkqCEKRFLEAYAUlQ1IEw5JclEM1pKhDGssZRTyoTUOmwdohXYejSG9OjjSmuptYHBEZGQsHGWEcHdqyqQO1gplQCFCCK4Tc1CgFZzMzW3cJHm0EWEm5VpsoiWSp6m6jGllJrNN06lWb3mE1PLXAsJqTsgSupb+Z+rpixJBIncXM1ylxGw1ppSjgh1a5AQAGgsDkmJiCJcMcDUy1RKmaqaA7MjqrsDgkiKXdQ6IALBjcERQyiYICI4kSckpGaFC/ciwkQNbtN1B+2ugIjaOqpaJzMNj5RERBC6OVMLLUjOiAARZhoEQGhVFaIC1LrrnIAZ4QDRYtXu7mEebo1R7eFuWmu4Q8Dq4oKZk6RpnLTWtjQqABHZAz2C+uF4pT/74M6Pfn73Z3fO10UtwrZQJjdtGI6PfLI9r29svPTFnD1GxJzl2vUrt269Uup0fHx8dnZeqkVgrcrcUDAzqwJgCx+bDegdRHq+X2pM9kaiggAgfLSbVknYSM/tv4gAAtz2QiP6fEv2Sc+BEIU4swggBTCgIGUiQUyEPMPPo+0VAplRCJiCKVpFgzsDok2KJQAdXCEMEIQxJUopy1aIZIAkeTLzIHD7Z//0H/2rv/jJszk6ixYtWrToaWoxoBctWrToudaa7t+yNwHsfFVe2t8XEiABakxGJIKEgJREUhLOiatWQGyLfNsWIiLMYuYheq1qZm0sAlufFxGQiIWRCIkIIXO6erD35jdu/eL2yTu3TxyxJaoIH/X9mfvFxcXVq1dERE03m03RYBJANKtEyNz6Bm2z2TAzAKgqM7fxv6mWaI1SRojhZg6PDPFtY7sbtNEJbhucIjzccV74OVcZpZxMq7lecvqe1/Hm100fcZ/hs7z4xfzB+fh37x1JObfNpmymOo3rC59qfS2tH8gZePzsTj0/K9LzyzieyFH1+uHto/X5Bbqfr0Z56Pfj3o0jXa/Wb713fv++ncvqnj6oZnfvX9y/PxHhnenknfMP3ru/eXBe9AvCFT7+iX++c+xpnZxfYer2Gb25Hnn6EVDNj87W3Xoaj1e1KCKaT8P+3iHnvsjpyere3XN3uMpe7pz2/fBwE0fnao6bgezU7qzw4YaIoaw0ndfNevXwol7goAN9cDatHqxC0t01/PrczsE7KPfWZQr0FiZc9PnVqLtxcXHxzjvvvfny4X6sX+31SrKBkHJq6+uxdQcCEgtJUmmqFgAAIABJREFU4pREErO0lQqMEFURqR/6LvfMXKuKcM7STEsMJ6QID4taJzcT5rb8v0yj1QpuVoupujsRMzeby0It5quiA4cjmDmyICeYeReoVc0dEVtQ+BEZHFHNSim571mSmzuYuWekZiUDMjGllFttn6TMzAgw1UqIOWUAcLeq2uWcc54Tpu5dzgBQam3XvqKlIe8BwFvjXE6IZM1aRQwEFBJPTEy4zb4iEEO4I8WMjQ7IOI/1mIWY5kNE2OKuZjb0QxJBAFV1C5a+9f3O7A8mpnAjj2ic6tmcRlRTgCCC1rTYKo5FRGsxVXMzM1Wtpd1veDuCwlyrAgYzOYSFNfSzqSKiMBOxlmKomMDm3C1agANJziRCwOdTvHf37Adv3/7F3dO7ZxUI5pQ1NDPVH2t7hPbj51mPPVhEZKb9/eH69WvXX7p+//7R0YOjs7NzpITIpY4sRsRq5tA+rmZnH6ABoOeFAAhb/vU2Du3o6IjckN/bW6yIlrunbTlha7ycUR3u2wqFT5qbI0QhEmIJoHCK4AAOEEQGgPBHnjgAIQmRMLWpi7aXwAB1VQMwxMAwZsydIDExS0opNYg5eoAFIMBk5ohj1NdfufLMDs2iRYsWLXqaWgzoRYsWLXqu9d3v/uvv/cv/PBSNEIBIsgKqmplqtVJNPZhT13XQ912Xc5drrUjUEM/urqp1Gt19HgiEtwJAZoloNMg2ALHqVqbRx42aSXeI3r3x2iuvvXyvw3cBMRDMZ8OaAB3A3Ver89Oz07Ozs9XFxcV6A7ABIARsGe0WfIbWc+iBCK1tqEXVWilSKUVVWw8hbEM5AOBbGOsMqQZoP2wLh1tMelfv7qp911ktVstXcZR+l/Wk+/zpCoCL9fT2O7/+n/+3v0bdeFVXd9MylVL18JfHV6+95+7H9+5N00SShoN7h4e/VNPz83MtBQNKrUB49Scf7u0NReuDo+PNen3wy5OD/fcsYr0e15s1Igz9h/3ecD7arz58WKp/mvP7W5m5v5Wh8eXzLp7pjp76xj+6wQCYSv3gw6N/85c/4PF0fXZSJk05l1q6vh/29kRktVofH52w0MHhg/2DDyXJZnV+dnamFgeHR1cPD48fPlidnwPi4eG9V35xp5RpXK/LNIGb/PzucOUdTN3FanXv7p2cO87D8breOT77LTHQ8cSM1+84iAMRiREj/GK9Kb8u//v/efbBGzf+43/397/z5s2rL1/rEzEYuDERMSO3bGPmJIgUAVMtAcjCra0PEVNKAFDKZOqlBZzHcdysc5Jw36wvXA0iJDEBRJiWEm4EwESMQAhu1apvucDRmgMBUSECIeWueq2lEEkAhtu0DTIzp0DYbC5E8t7efhKpUKtuMpIkMfIhMRP1wwCApWg7M/f29opWNRORnHNKya1VGkAjXrXcagCoKs59fUBESaRoMTckmi92AITzmiF3N3dqTYosc7GcNY5FILXrpppaRHRdBwDm3tY0IXIrMCREIAJEtdoeVUoJPKZxojAkyDLfNkSEmRZVnHnQ4RFmXkpl4pSkagUIJoIIUyulNL5Ww5uUUhERWyAXMALMDBEa55qF+6FrsWhVm6bJww/3DluWnJEacDjnjlgkdRpYgSh1eTiQvPfDv/je9/72F2/fPjsrpgDm6O22BBngUVj3eccM/QYRYd93L7/88vWXrnfDcHxycu/e/fOLVe4G4lSKIU5E5A39PFM7dh8+8/wOXXLgY5t+bvMryA1Bo+3V/sjdV7OkZwPaHdzxUQHhPLf06LFud9sA0ELADmRA4HOyGj0IghGYgImQhCVlmc9KADULM6tazaq6mYrQ0KVhr98buqHPjV4OEKpVrQYAECN3JawCunlkMXv608uLFi1atOhZaDGgFy1atOj5V3BfQZNH5W4fuvX69GS9WtVS2xpZIg/TWiYOQcRGlGxDCXczrVXV3QKgxVsioqoiEuFuoSVi63dDoNawTghMb7z68us3r13d54dTFAXCtsazdfpgAJj5NE0Xq5W5IzTGJRIxAkNEG/ECQK11Hti4q84ZZ2Zug+qWem7LgRubsv2wDYp27vOOadhG721w2x68AxAzscDc574bgiIA7BpznvYo9OkyhV90/XZp3PU4vXf73r37xxEWES106mbmQHy3xRW9JfdxV8MV7m2t8VyGSfg+Igagm3sA4X2cVxDPx5+wwWpQLfxTDtFv6xt+rJf9sam759+RfCqJ7C/yNC8/gHk7U6m37xz9m7/8YehYp8ksmEVNGxsAANx9GpUZc5dEkoeHWVE1c+YPckqqqqoQkJJ03bsQ4W4t0KduLAlZ3KOUEZABqTqMtRVcfr5nvay6eCxvaRFjqXePa1g19/snmz/59uv/8Fuvv3TY94IQjhjE1NrzEFFrrbVorUAQSmrayswmAHcfNxt3R4eGdAZ3Y0IMdEd3cHdXh4BwrdXcW1MZEYKHmrp71+d2oeFOuDFeGkJCpPlqRAyA7p4HAwARkZSQaJomIs65yzm5+3DlsO86EWmnChIKcwTkzgCAmUSETDyirQFymD/gCIEJMHzG6UZ4LYiIwabGROSiZVLTGYKxbf01RYDAAAF0N6sBxG3y1dRie7lsl/jGJEE3MyuliAixEPEW70uAGBCmZqbm3nUdRGw2bZYaStoAQNuIutZaAVvEGk1N1T0wSYKAqUwRTsTbeWxnFkYOxGChDG3au09dq627jCRm5pRFtZIpSdrbGxCRSLjNUQMhAISLCBBXD9m/gt3+0dnqVw/Ob9/94Ac///AX987OpjoG1BZ6fgTMhvkk3J6R8Uwu/U9d8ydJY2aw8M1bN/cPDlfr6d6Dk4enF4Fkge7hc4vzx3zitqpAACJEn+99HpEz5ruliFB3ayQYfcyA3lLOYrdizqIhMy5jPR49/0dGPzIgB6AFeqA3GgphhAhnoo6py6nLKScRJiZ081EdwtzUTcGtzaxkyTlL3+W+y50kIQZwcHcIIiBCYkQR7PJKbXI0iGRRd9H+RYsWLVr0fGsxoBctWrToeReJuwuDT1Oh/cNIfTVYb6Y6TUPf9ym3jHFxJ63IREStKJCZ2iJYm2ve3FS3jrC6x46p18a6EECEREgiToSEt25c/cbNqzevd6sH01qdEGO2f2HrQYeqrlYriEgiHrUNnEXm4e4OptE6hZolbWYirXh9Bncyc4vkzPDKbWNSewUuN+rMoE/31tUecyQHmZmYkSXcYC6HfzQ+e5Ye9KIn9ekvSwSU6q2m8qN/aAbwZN/Rb2pAetJeeNIHjCe++Ig+n3n6sX91eU7i+beed/qCcOov/kw/ugWP2FR9987xpZ9VAAB4/PTQgKkAfGTpgwLoo+9KhVXZ7mY7oQV1u8Entvn5hS/acX/6aov2d9+ODrdPNvdOfnV0srlY297B9a4/HIYevEAoQLiBVQ3TadyM4xrCAwMoSp3clABMTVVNq1XT6hEuIn3f1eJE1Pd9AHrMJlnMFF10gAhEx/BQQwDa6/ZZ2My7lEUEmYgZid2jRXe36znmCw0zszAxxxZbnLtMhIemNBMedlO6Ye7Ec4GBhxMDIRNhVS2lNI9YmAICzbXUFliu0xQBROjmCEBErachIlLOOaVt8NmkdQIS1VLVlOYdxVzGi7tr5XzujYillHHcNIIBkbQLKDO3B+zuZmpmfd8D4lgKzmY6tbldIvTwqg0/gohcq6mGcAYGnEPNja1hHs7ClEQkBYIgAEaZChMfHBy2R0ZEbUIZ25MHmKbRTAmh6zoRWW9GRMwpZckEGGa5T4F4NpX+6tXoD4+Pzv+/X97+6+//9Pb9i5N1NYIaYI+5zLMvuyMix8ddIZ7Kaf70NrU78QDafRWEpPTKrZtdPxwfnx09OD1fjSw5kDwA2n0Rwg7TvN0IeLibI7q3cgykdqTn4DNSuxNqt2HNeoZLy84uP6vtdqMl32fg2ce5+ttQNUogmaM7hxMAowtSxzSk1CUeutx3WSRFuLmWaqrVrRHhTAj2+zR0fZ+567Y+dVtJ4R7gHIBITCKJqetUpJoaYqQqm/zf/q9/9fQOx6JFixYteoZaDOhFixYtet71T77733z/f/yvJqHNVE7XI096cHCly3l9cY4eEFCmEuGByCmxMAkjETOnlHMG9+jDVbXU2gAc5rbZTOM4lVKmaZqxywDhSoSExMSBCbjHHq7t599/89bR+t7perWNBl5mpGIp5fTk5PDwMKW0ZTjTnD8lYuad+7zL4rT4cxvzmNku7ExEiCSSUkoiAgBtdL1zn3GrRvZoC3tb15Agt8BjGScHay3yX9oxWgQAL4Id/1liy18bfY5A7icn+p//4/vpimduEH+mjX8dw9JPTvOgb40yRXr/6Kz++O9PT0//nT/85p9+55sDeyYX9DADNwIIrxAmiTxMrXBKSFCtggdFEIIkzsJtuQ4Rh4WZjeMY7gCRUp4BT6yAJF3XoNJEFBCI2A8DIJhao8k2ljEA1trmZdFMt/OmAQDuZpNGBCA0yrFsxCNqKS1a3Wr+Wq2bmdVawwMJU0rbq9ZM3kAAAJwQolYwI4hWDjx704DCEuGNYtGyzL7ZlHEiwgbINSa6FGh1xMav8Ah3K2ZJEgDWOnuLhNgiyT7zOXAqRc1SkpaCNTNh3tvbCwB1j0DJiZnMzcPBPUuHwOAhDcIrKWlYDfNIKfV9Lyl5eNsaEUrOEe7hxERMSDBNEwRwYoBoNRPUjFAkM6ulEjMgQpiqmTkSI5I5nK/WZSzjZnPlpavDlav5yvV37xz99N0f//Ctd/7+Vw/eu3uxKlYCwMEbl/oRnTgun4GfCl36ytVCyQAIgQ2m4e6Hh8ONG9evv/SSevz6zr2L1UY1oJ0KLQLQ7m7iiVucLUMDLi8gozZbMd+AxXavO0r2bonZYw/s0UsXEduSw497LQkgI2bADJgAOpGOORNl4S6lIaUuSSKCiHGqth7N1UxLmSKcBZOklHJizDmlLEgRbm7gSIhEgERAxCwsiSUxZ8aULRCQAGK4f2hv/PqpHY9FixYtWvSMtRjQixYtWvQiiOgKwIU6X6yvdZIYCcFKsVrDbI49zYPKMDdiRoCIYBYWRHcW6fteTRvymSXl3G15FxYtOWOtoT7c1cMDnUMOO/n9N177+w/O7jxc1cdKaOZxda16cXFx5cqVfhhIFAAiwswbZ2PbVzRjnYkYoMXNuIVrdr/Whs1dR+0XGqCDtijMFtXBbUVhs7MbqHC7cDQkpZxzLQX8+R50ft30HEY+P8F2+Mg/PfVH/ly9Gp/bfnnOfZsvqK/+GH1NX9yPLjRpvXBtQf7pppRa1uPmdLV5eHz2xo39m4f9tSFxKIUnBqJA8jBwcHNDAgjSqjODp/EskEgEAN08px4APIJbYZ9ITimlpGYAQCJEvLsAESKLuHl1Jwhwd7NADAjXed3NVEq4ExGAt+Rliz6bu5m6OQtHgJm28rRmQAMCkYSHqjZKrpcKAN7KcudaX2wpadOZNkCEsWNAE6tVd6+1NnMcINRh63BHRKQQRAxvdXHBIs1ndHfVUDWgRIjq83XZARCZkxBsL8PuTAQNVhBAbcY6Zw8gc3RCSZwTQetFNJBEiF3K25eRU0fh5G45577rVbUZ0ETIRJyk2fTUllQRMIB7EFF7CZt16gDj1BDZrmruFm4tFg3UENlk1dTciFW6kdJ6rT/+xYf/zw/e+vnte/dOp7MJrD3B7fs4Pu4k/JhvnmvFbp3WlStXbt68ube3//Dk9N69+6UoN8LY1qee2wUfZ47A1kOe+zEA2zR8QDzGzbiENdt9tZvjv7St1mbpbXEBREOob/9tvv0LBGDEjrhH6ZAyQC8y5JSIEnMSQkLzsHCr1WpVrREK6ATBgilRl7lLnBhzJhEgAMRAbMCNAAgmkiS5SykJJwZGSHk9lQAIc/iz/5vf/dbTPRKLFi1atOjZaTGgFy1atOgFUAcwajW181jduPKKl43aPLAIAE4shEjUxo1ugdRcZiEiJnazlNL+wcFqva5aiWgY9lue2NxUtU5TLVVVTVWr1lpc3bWanQ2JvvXGa9f2f5UZNtqAFxFt9IMAAC2DxiL7+/tZrdaqqoiOSMzsHkS4W/bbumIQoTnLqtpQGw3BAQAtO9aghLGtZP9YBIf7o+XPDcVBwpKEiAw+GudZ9Iz11Tt6T+ize9CfT7vFyL/pn150fb096EXPSk/ibwLCQwPBDVYn48PzX7337u1//4/e+JNv3hxu3ejJhV0AG/i9lBKEJCnc3UENkZCIkdt/JCm7h5W6d3goKZVShmHou87cc0p933uEa9VpahYyQCOCYFTTUss0bQEU1i4qu4vROI4I0OXsbrG12yJiM40RQEQiDVJMWtXUGqKaiFCCkBIiMbt7maZ5ltQdiYgxPMysaIU5t9omej3CJaVEMk6TexAJYyJkREQCdy+lzP2F3FYm+Wba1Fq7ASUJM1dzNVBDDmJiRWNiJAoA5IbtYCQy9z5nb0QG84ggZiYCImFBh4oFkmDOQ983eHSEtXnriF13cc6SCbGRu6bN6KbY3GciABBERURqEd0g4ga/nsy8VosAADN7cPSwVhXJ0zSp1nBnYWY2QJ6ZYKnb27ty5Vq+dv3C4Ge37/zNTz74tz96f+UwBShsfefYmbDP29Xnsyq28OoGDGnLBa5fe+nVW99IKa/X49HRw4jo+k44tRn3nX18ib9xaWvbVPV2nr6l5OfodPs1ori8BUQ093j8lqnNugCEI8CcgN6FoHfuczBgAuoo9SQDUALoJXUpMwEBuPumqrurh1V1VQgVgZxwf3/oO0kMnVASYoTEQWhEyIwiKImIINxYuOu473PqEolUd6W0HjcGTg76sz+SP3zr2RycRYsWLVr09LUY0IsWLVr0AuhPvvvnf/k//JfM4ubrabLNVM7PrWxcK4LnLsu2fI+IhNncXHW9Xq/X64hopfPnZ+dqCgiSUt8NOXcQQSyJuc/d7PU2C7oWU1f1Ur3bp7x/9c3Xb7x7dHx2tN4NUmKHDowIj1LKOI7mUbWa2m5w1Bgal4AbvktAu8/Q55Z3ji0wugW5AVpGrW0KmbnW2rJXiDSvPvaY/wuzlrFCJBEy87DFg170LPU72D73mwAdL5z788I94BdbWzLy/Im8drg/+U/ePdJNLeP0xivXbl0/2OtzToDsEh0KsyQUAaKYA7zMPCdxmxPXyvHCHQGmcdRaU06lTCcnJwGB4eBmatGmPAkR0arWUmqpxNQKDJoXTMRqZqrNrgU3LVNVjQgRIUTXAkhIsl5dQEBKmZliburDCGQKRzezBhJvZI824eoWboFEDc2Rc0cs85oehC5nADD3/f0DImJhCHC3UmrXdSmncRzbSqYuZ0SotQ77hxDR9b0IA8B6szFVAOj6HgE34yallCSZ25bcO79+zXBn5hYJ37rzkHIOpP3qtH2JAyJiJkSbWd8PRFhKcfPRNsJSa4GW6HZzdwjwVnjIJMJqVU1NDRGYiEXW6/VUJiZxd1MLiwb4HfoeoEdsfF/uhqHrh9T1QVmG/f7K9e/97U+//9NfvvXug/d+/XB00KCYZzTmM+tLP5efgeapjpmbwUwv3Xjp5ZuvnJ9fPDh6cHZ2WooFkshlfxkQkbdry3aySwXOLSX96CM7wmPmD/nlW6Mtl+OyAY27GfxH3Y4Buy9g/gIBGCAhCgRDEAEzq9Wz840wMQKGm5u39zASC6cknWCXqEuUGBJjEs7CiaB9wUzMJIgATkTD3pCTpMSt0aSoBksJLRBunsN//Hb9n/7lMzksixYtWrToWWgxoBctWrToxZATFabDaVqtxswSJEgEiH4p/bNdkRmubm7k4W6q5hFIWMcChMwUaugQ6tuBDLIwtxpCRCFKzO5hHmWqA3XDle7Nb7z8yvv3P3i4UfPHGdAAABExbjbrfi2pU1WtSiyE4O61asScdEbE5kcjIvOM1NjGc2Z2YfuF3Q/bCJ+ImGkXW2v5ne2vQBsaRUTjRwuLkfrjlWK/C+7gos+lL56ee55NkOXEf1LP8/H6mqs5bSXgXONXD1emVsI2BsbC3cB9HjpMaCTMOSEhEAYiACFgI9k2tG2EY3gp1dRmDxQgd7nWul6vAYAQBNFMwYOYASHcy1TcvDnO0JpsZ1YBtTdKzh0RmbtahAOJIHIgECdmSinXau6BxJISMZspIhFxktQ2GNvGXVVTNZLUjMKtu4i565llS66gnFOtddyMKTXfWMxMqwZgyinnrvEWJCVhBgAW7rogoq7r29WzZa4BoPX6ImHuupRSrXWmdUC01UjEBAHMjIQI2ABc0frqEIQRAMDNzGImkLip1loFERHHzaYlvoU5PNwMAcyt1urmqlpr7brc5TSVYqbuQQgsknOexlJKZXZV06qpy8KJmZuziBiIyCLD/l437HG/vzZaKR4dr7//1q/+4vtvv3d3NVY3AAXwR22pCEBfi4+4Xao5JPH+/v7V69f29w/uvfvew4fH69U6gJEYoAX2d9Y7CvMORwYAgGhmHr7LP8P8fkFokI2PobQHPIGSxvkRAQKCO7Tc9ZyAnrPPu7y2ICVEAUQIhzAw96q1iCFhUIS7E0CSnBLlzEOXusx9IkYXjsSUiIWICRJzTkmaB03obsLUdR0ReAC4W7i6A6b1NCmAIvzX/8v3/+wPX3vGR2fRokWLFj1NLQb0okWLFr0YUqauVkVY13r16rWrQ9b1yTSuap12Cy6jxYs8SqkBsJcSsbRK+5Z/EWQC8qIXq1Nzb6YwAEhKLMxtCApIxEzMSF1OlIe9dPDNb9x6/ebdv/vF3YDHnV0AAAiA1WolOV9/qY+IqjUBBW6X+3pLmRERtUFv22kbcgOAme3qCmutOzO6LXluLYVElHM24509DQCIKMIRFBDk3FZST5tSsQIQbFHQX4MR6qKnqp3pHI9/+0X0qVv4Mk/Dy8/u6epr8Gb6BHbKomejaKZVYxNjAFSI44DpfDr6+dH9VX2wqZb2vt3v76c9gsoJOSWgsDC1GqZhEebgHm4WVmstpXrMIKp2MC/CTbWqmjkRpiQYwczdMFjVaRpLqZJkbxgiolbdlA1TJhI367o87A1d7tx93GwCOQ394ZXDWmupdeiGlFJOKQ2HACAiucsi0rzsRppqxW8NeZxzXl2spqnklFgYCbX1E26dQQJMKRGRai3TWGshAmFEYEIUoQGyu43rVUAQkSuM04jbOl9CQAwz1VqHrouAqdZG1hDhZuGpBmAgBAJGeC1KhABQSlVVN0OkcDczJAwPrTpfqwGq1lqLCDMxEW2OH9Zax80m5y7nrv2+mwVEVd2Mo6oGQNd3Dj7VUqZCxF2XVc3CAQM5pUzeqNiAXTf0fS+cct8xS4R3Xc45EQHm3lJ/cV5/8t6dv/p/3/rhT9795Yeryd0AHMFx55U295kuG6MvrKghzt005/TqqzevHF5xj6OjByfHp16VsuAMMWuv4AyHMdWGzHazAGAinyEdOwoHzH7yLmTd/rf78Gtmc8sUbDPPzaem+ZbSwg18Z0DP5A3YthQKkRATkSMWt2JKAJRYw8iDwwkjEe9lHrrU93mv7/osSShcEUIYGQECzCwE2l1ikpSTAHg70TfTaFpzSkBogFZtXYo5mdE/+w/+4b/667e/pKO0aNGiRYuehhYDetGiRYteDP0n3/3zf/vf/xeRsJgW00S02qxdK0AbXgQEttW1YdAKkabN2AqYgHD2bZGaKxzuYO5gwswiFOBV62QsxCII5OAAbubCyhneePXmt75x61p++8Rt9EfYQoB55ehms+m6nl8mQmpEjvaPZt4GP61RcJe1aU50rbWU0tYFt2FVg288KnAH2PGg2wOfozxzejrcZ0YHELqHmbOwSNJStyusFy36iPATv/0aaOexfu7zH7e+/OUtXHbqX7h31u8IJuVp6ena9Je3hgHggBVw7VHd8MFqsjunq+no26//8e+9erjHw5Byr6VsPCozhnqYoUODR5Q6NQDzXH8n3K4mrYRwQHQzJExJwg0RU9epEgnuHeznlHLX1Vrc/ODqYeJOKLlDQw831HHOuTErJKecu8GdmBAJESTntlNExAaDaI29bU4UgYnDfV1rKcXNlDDAiUBrdXds/XAACGi1AKJq1VIIw7SWiPD5Wlm1EhI3KrbpWCaIAEBlImJkGqfRzNxsM66ZGBDVrJUM4wqZCXEGWzfyBjxiLUD7YZIUAN4u0BE4G4+IiF6K10LUI4RWgwBBvHJ4AIjhUaeJRfq9npnUPPUZIhCRRNorkXPfnMQ2l0zMIkxIatrqI5JITqnLfdd1SFSKVtWL1RSEm7NyPD783k/f/9E7H/7s/ft3j89Hm93n+MhnT8DT+KB7HhSNYQIRwzC88cYbOeeTk9Pj49PNZgQUSQmJzVrMGZCa7Q647cMAREKIdvDoMft53kEQtD/e7W/7L9vsdTz6/faPrX7DPcLn27145D7vhAgEAGHm4OERxgSCRHMttifmPqe9IfdJOiFp+DRzs4rhYRDMIpxESASZA9Dc1RQgwEMt3C0AVGsQGeep2qRQXWmCN69deQaHY9GiRYsWPUMtBvSiRYsWvTBCJz7ncdBpWnVdv96MACpMAEYACJREmBhwXlNZagUilgQB4AAeYWaODdpIiOAOzIQIEWY6lUmSiEfwHJIxB8eapNy6cf1br71y82pXzKfpiQx0QJnKNI5mjoTEXKu2ccpumbOZmTkz7WDQrV1wRhYSuequxB13Y+XZQcZHtI22wwAicA9VJ5whlw1YmUQsp1qSqS/+8xfWiz62/1R9jfkb8HkPH17629+0hRfxxHgRH/NXpaeyLGC3rTmKGYDb+lp0gAJQAGw1XWymO0fHF+tpM9bXb155+aX9K1e6aXOOoPtDF1pdjQNTSiLSqMPEjIjM0nW51mpmfd/nnJsfjQgi4qYBTsKqKbv3XZdSIuYyTQHQ5T5xZmT3GeJUSo0IIhQRQCxaW6ttW7tTVWeZ6fzaAAAgAElEQVTkAeIMSPb5UtiSqRGRJAVErdXUIsItESGA11pbjSHOaVNoM6nWKBkRVl2RtHKbba21iiTICQC0aikTAESAh0sSpAZ0dogwM2buul5NawuAb5HQAKCqZSoe0UoCAZAYVdXMVaw1+oYbRBAiEzEiEWASIexyDghwJ+aU0jAMRXWcpmrIifu9TlICgN56JkZEj5hKUbWh30MkUwMERAjAruvaYiYiYiKrlYn6lIjQ3FV1vR5XU50c7p6t37nz8P/4m7d+9usHZwUMwABidvsBAPCRkf71eS+3isCc5fDw8PXXX0eiB0cPT45PxqmSJGZBJDPdgjXmzzFEbPdQbfWYe8zs5y1/47HtX5I/9l3b1KWXE+dAtJtvV5vFFvr80de8cVvcAMMxAjAiEMAJsaGc+y7vdXnoc2aWdtPZuNBhCAEBSMDILELMAeDuGh6O2/eJEyEhmJsHGuKqTEps4QjM6k/1OCxatGjRomeuxYBetGjRohdGVLh2G8bQMkHOLEmrFq1uFTwwsO86YaGAJJJSSqXQ3O8HZgY15sSWasvJtOFFW5BrZuo6jgGIzMwsLFnSoFE25WSvO3z95rU/+OarF3r35P75Yw8rIMAhoFY9PTvdG/YODw8367WZb0dBiEjQanDcmpWMCMyJmHY0zAas3I6wEFpQxixxIsKWfYYtNtrnsh3q+34evuG8p5QyBIT5eq3uT/JCFi2Cz2BefCrF4rPYc086nk/T13tm+ozOzvP/RJ7U8/KYnz8v/Nlm29uimbYPmvcyk2VHAHUYK/zw3fv3Ttb/+A9e/eNvv/advVsp7+2lONzLVkctBQJZkkiKJIDQFs0wUT8MfURAdLljYUKsWhBAUjJTD0MkCQeALmVmIcLcde26hR6uVUudHTp3d7fqbuzu4zgmSc05bSyOZqF2XefuZjpNEzM3mEZzk+va3T3Am5e9t7cHGKa11krEXe49MAKgFfi5E0JVLdMUEUSUUiYmQHT3UqZYz/OvCFCtllrLVCRJw4EIM0RcnJ9HRNd1MadYuaqaaZnKDLkKCHOz6IchpwwIE0yTFw9ILMMweFiYuxkTCXFKqeu7lPK42XhLf7fQejgRZMF8OACAopsVFun2+u2ksu2lPQRMkiLAqqkpAIgIExFCSqlqncaJEcxiNW5OTs5W67Gah/QTpF+fbH78yw9/+Pb7t8/XFwogENZOzWi1eM19xnlqusWpL5+0+Py8wX8bzdHmK1cPbt56+caN63fuHd25e+f09MxU09y63PAUWwN6RnvPK9uYGQEN57ud3QKyL7ICLCLcNcIiDPyjnBPcvdbz0jRnAEJkRCFMxEIwSDrs+iFLuytFCAd30xajzjmJECNIkiyJU/KAUhTDEYAIiZAJRURrdbckhCQRYE7F3U977PWf/19/8wVe9kWLFi1a9BVoMaAXLVq06IXRP/lP//zt/+4/O9qPql4sDq6+NK1PpmmN0TAXWKtaVWqV4wCmysQhgYjzIlnibRsSzUsnISBm9B7Y3FSDbSSuaj4FmkPtJR8O6R/83q13753T/fPLy2F3CzprracnJznng2Eo07SN4cwB5W2URtowpq0bRaJWKtSiWARAPA+z2ngeEblltMHaMGzeZUBrLmrfIkJs/5aRcoT33TStG6Fk0TPTizja/9J0OUf8leg5czgXbfWVnxnw+Fv3S3sY8ch9bpeNCIBANsQp4uGo5eisEq5VN3X61jdudK9coa7nlHOvCNDmRQMBCYm4TBMAdH1HSK3rr7UJBgrE9kLXCgxZiNADwCyCzB3AEVDHolNx1XaRAoi2jCYmaPwKV61EtdbNOG42a0JKKZlWM2uzm6a1TCMze4SbqSpASBIzjYjNJgihJZoB0Kpt4cXYIsySkpmbz1aquambBwAEUgtMQzSrmjmn7YkTsGtN6PseAHKXvdXwcvJWvBDBzCLS5b79VddlkQQI/TCoWWN2iYgkRgirioCECNEq41Jjd7S9BIC5h07glPvscz/w1uXEluZWQmKShuKepgIAhAhhk5mbE2Gb8K6lWFVXLxrVQIGPT1cfnmzevn3689sP3n9wtgqoOxrxVjuAy6UfPjm9By/gVQkRARlffvnGzZsvk/DFxerBg4fTWNyDZ/5Yw8MQbqnNsKsVRDRznKd0YkvV2HHLPubN/fgL2PAau5c1mr3t4R4znmX3a3Hps2tr9rdZJCAkJmSAzNLnlAh7kS5lYUJqILVAaJWigEicWISZkIgCoWo1CIygAKbtHSkTYQsocAAisZoHURTHvRLr/MyOyKJFixYtelZaDOhFixYtepE0FPqP7h58/x+sx1JefenGmiDcAinI3L2UUtUIwMzMHSNEUp6L5jFaroRZRCIQAUXYPdrg1sNEZ3Cze5i7WtRaHSzQZFoPKX7/zVev/+xDIdjBLS4PblTr2enJtWtXma7u+I+NjkFEzSJPKbdBtara7EnP2yBuj46ZGQndvdkJ27XD88LSxvTYIgbBTHHLgGbiufEdOEWen/WjAdgLET59nvVk3OxZ7OI5MeV+009+2y3A40/qSd/vi7yMX875jC+ss/O11afm8z/hr+avERG+Akz+9sLxaEULEiMQYFTXs2pv3X54slodnx47/eP+8HA4SEPOnUBiFEKmBjhGRFgTmFlqXXkI7u2S4hThHtV0i2YOEY5o5A1koqIa4cI0XqzLZoMBKYkkbsFkU63V3AOJVB0gVPVidbG6uOi7vk3Y1lIAoh+GWkqphZibJxtuLEyJScjdS52YWUgA0c1HHREZgQCosac4IRJzynO+FaCqmjsgZpbcZQSotepUhm6QJGamquGxzUBz7jpmSimrKs5XWIptywIApC3DYZs/n1O0EaCqWnV/fxBhq9qoC2WazC2K0+NXXmLSUIcQSQDRPHs311IaxKvUyshBEgbjOK7X65yzCGOBzWbTaiFEGIlOTs6nsUZQf3gNu/3i9P7xyY9+fvtv33nwcFMnBAVwAHPAePyk3VZO/uaT9oX8jEIiEXnl5is3Xr5Rajk5Ozs+PjW1QHKPxmM2M0TfPUFEcA8kJCKrGgBM1Hov2lQ9IjbK2cfs7tFc/rbOY16NANhC5jP9+ZErffl/zXpukWcCoAhGYiIhZMQsaUhdYso0f8K4QbgTBjMQITPN7ZZESBgIGuaq5MGAQtTO0dabbWYpMzGbKqCoT25mAqHxL/7q+8/sgCxatGjRomelxYBetGjRohdJbx7nn7w6Tu7nm/KyYwCDUeZsUSedmFiyMFIpBUyZSZiBaD1OLco0TgURmduoBrsuIxIgMgQySU4iiYja2BsAS7WqbgFJ/Mp++vbvvfr6rcOXDuXhhY0WtgUybgM57gZWNdy6rltv1uvNuu96xLSrEFStbQRlptpcckJEVFUmRsJaa8s1t9JEDw8WQlRVmPeyZUFiM6CtmdwYFDNVOiIcwLu+d/dpHHd/sWRCn4aetaH/FLf5sZt6Hs6Bz/IYXkgnZdEna8dChq/oRMQdEQkAAhy+7EdyaV+zDepuAW4ABOGIBPFgXev7Z8frv3v7vbt/+kdvvnnz2q3r+1f3JJMLGIEiODhotYDQSaLFlbWEGyDklCOoVGvlAWbm0bC3Eu0yAe16ZLVMoZpSTh5UdZwmAEgphaE7WFEiYpGu3z+QLvUHwzAws7lx7iMCkPLQd/uYujyXKLR6va5TVXcTkZYnnWdikd3BzGu17XIdjHBzo5lS5SknIlbTdqVjYgBwdxZu1CxmJsKWv8ZLSo0f4o6EhGitmTgC2mInjFKKmiEhixBxLbUBqM/OKyFQQOtnCAfVWlWhAbvMmhuobs0xLJtN1Wq19MMeBEzj6A3UACAkwpmJ6zhOF2vszQjNCgAKAgSQGSG8dP16yGA8vH//9Je/uPvWux/efnhx93RzPNkYs/vsj+4rHjtjZvDDUzppP86f/YwfvJ+w/4/8Ez7xxe535t/MWQ6vXrn+0rXUpTt3P7x//975xUUAEs08lm2N5KMtN5ALtPppIoxHTZiIly/NiAjh24pJQEBoaQAAwIg2GQEtkoANy9x45vG4Bz0/g4ZAIYSOZUg5eyQAQeY2OYRARO3uzYAYI4CAkChh+PxQ54kWU60R1uXMIuHhbohAnFmYJTEzE8j/z977/Mh1ZXl+33POvfdFRP7iD4mkqCqpStXdNZgBXIAx3vRutv4DGvDGwBgGZmcM7NXs+g8YoAEDYy8GA4/hAbyYvWEvDDQw9kw34EFPu9vTXVVdKkkliaRIJpOZGRHv3XvPOV7cF5HJJEVRKpJist9HgpQMRrx48d7NeO9+7/d8DwNAqaUvWWLXq1Yg97XMr7zYaZqYmJiYeLOYBOiJiYmJywT94R/+yb/4J2whQ0+WA1TcaayV9M1UrdmciYJwaw20/Zsx+IKo2aPMTISJhWubOrg7QggOCkTMEsyZyQGQ74QY57s//sGNH966c/rpYdZqzYaDMynSzYZ+vV4t03zBxFq1SgVaE0Jzbz0JW3ChWuslBXG4qoKdeMzHxKa+1B0MMqBNrs6rz5ugwzEvmrav2Lh+UkqmOgxDy43c7OWboD9eLp5z0C6jqfx7HwnTCPxbyrZ6fdNJ7SVv+Tmb3ITxg0A8BiOgpS359/ZbPL7pJkqg9ThjJj8tWJfyeP3g8HR9tC4/fHf/h+/ufXBr95392f48iGdxFYeq+fhZzGod+hXgQVhTB3DOJiECXGuuqg6azRJTqGYi5HA3hJAopNSl5vYNTsw8n89NvXmNY0xd14UYzGxeNaUIRy55NAUTiQQJwsK1lpiHlFIIgZk5F3Obzzp3a30ChYVZVF3VY6lBAouYqnlL8yAzrbXO5ouUUt/37ZL35JWONksXHoR9g1rryzhqhgCc2cxKraUUcxcRdx+GIZfi7iEGkZCH3GI0mCAgBgURYTbzYRjyMIzB1qYigYjUVEIgpnXfay2AsxMTaSlmCrgIm9VcLEjwquzQnI0B9zTrmGW1XoNjjDOV2Ummrx6d/OUn9//qk3u/+OzOUa9rhYIM1FpCtgFybvH4iZHzir9Dv/HX4Rvf/xnZIU+WENF5DXqxWNy+/d7BwYG7379///jx41pKCB2JjGUKF8zIm/CLTYzNM/b/bDSA0aTnMUfj7H3JxwSVbbsOYFy32KjPz5b6GRSJZxLEVdwFY+0ZUQtDr+RsgDFVUwcJQYgIZE5QNxi8EowJSBREHKDAgSEi3CodmIiaFm4Gh4TBcnVSo/vv/r3F8qtvOgUTExMTE28ikwA9MTExcckgl5BD363uHx3uhEiOYRjMKxy1VLgjRqbmcmJVM7UUO2IS5iZAMzOVUkrJeWgJGWNTP2iadSEmZkkxhRDMLUhIKalqinywu/+7P/rBr7589Dd3Tr2v1DIjx8BKAHDH6fJUYrjRzUSEmUsptVZialmC29TmVoDMzGPAoZm5k9HG/jxqzS3J+nySxvg4kZkxc4yxPdJmy+3B9nJJSTe+6e9bc7xEXMjZuPDg+T/6U898bTLWd0sgeOZGXi5fp+U9PfYunXA/8bIY9cRn2i+f/7LvNuJpE7jRBGh6I74KnzH+3UlBCiY4E6ppPlx+dfjxXqT3rs3+07978+/+zvs/+cGNhJpgiVFrVVW4JxGC9+ssDJl1eSjmVNXnkiQE1SoMkXRl/0qIs2rOoclkBTAWijGamaoSU4rdbDbPeSilmNrO7u5sPuv7vtZqam6mpiFFEQ4hzmazFvQ0DEOpOc5SCMEdOWcnMBELu1MLrFKzogYnAscQWYQIqt5Ce2vVnHMehrbNYRiIWERqVTN1txBaPJWcnp6WUhaLRfNBD8OQS24VQsLSdZ2ZtFXe9Xq9XC67bsbMZlpKyTnnXEQkBCmlqFZT21ksggRX61IKIn0/DH2fc27NFUFYLCSEEDgAqLX2qzURdV1nasSUYnQPBIoxDsOQy+DmBFrMu75fwWk+39nZ3Teih8fLWdctdq4dLfNfffblv/0PP//FneXd4zyYZ6Bu0rEBAAqc995u1ipe+bB8RdCTA/7i9Wtvb+8nP/nJ7t7+er16cP/hej20eG4wtxqF0cx+9vr2m0xw2CaMm5g3MRo0dgZUcwexswhtGjuPxQAAgNEI7a0p9eZtzFzVzZ+5StZOkoxB5k7mMHdS+BiXYo6i4CBOMIOaERBAXUqSgtZarLpWhoZAsy6lGGepg5sECoGtVneoGwPqbpoBUAhpvii5KmCBrh//5uH+D1/OmZmYmJiYeL1MAvTExMTEJUM05NgHsiHbPMTZbJa1hxEDzDBzU3UiB5nXNk1hOMzraIeBqhIQQjB3YQkx1FIVFea1r5qVRQZfN/tVSqnrZiCnvgwZV3dnP7797vV5WC6xVEB9O0Fq2kYehvVqLSKLRXJv0RkuImZm5ucF6DYBiyEwCxOp6eYJ23pTd7iNyvX48VW19V/aStjNKbZNnT4Trx0xxtR1NQ8tKvrSTl+/F75OIb1QUHz+oL5+JfoN5BsPwvMPzku3o74BYuMr5DJ68M8YpegXU6IvftTNiX3+539q7chH9crf1GHh7oQm2g5AcdfiejTUv77/aOkPHg8f3Di4fW1vZ2+Pcs81u2lMKYaQFgfkJuS1GkucLXaIWl/BzCwhpJTmakRFiYMIRYqbfIvKRMxiZqpl6M3dmRzkWnPu3bVYLbUthZppLUyRDJrdiNw9l9yuaO5mZjoMrWGcZVbVWkrXdeaeh8HMhaRLszJo1TpKhW5mxuazSKVf6rByVWJxFyu5NQMsa2vFPSISiPrTk1JyKZm4pWizw7XW4+WSiJlFQtBSULXYOgSJMam5OOYhSBAR6URUtWoNwkJAEMBKVbVCgbrQdaljYjUlJnXVorlqqUYpCQsFMaCqaT/M5jMROVkPtVZXUrPmqt7f21ez0+V6ceX6bPdK1+Ork/Vf/vUXf/3JVx/fOfzN/dOjVe3NC2BgAp27zl8cEwD8Mv+mfx1ECEn2DhY3br6jqo8OHx8entRqMXUiAgBwBjmBIOdehtZ1E0C7rWsh3aUUM2MmIoaLtS2MdmkACCyAbG6wQJsvHmZiBlpWx3gH9qyvBx+ldAaxA2ZMFIQZxEIt3zkQ4pjl4lpNGMJEzKXUmrN7jVHm3SxGioGDMMC1KtzUUKvDbXRLkCSRWTdXd+PgHIzdqg4r/eTozv/+f/zJqzkhExMTExOvlkmAnpiYmLhk/P1/9If/5n/6J1UjISsszudaVl6dYGKCCrcmBZO5E4FHTdaaYosWKLlxxBCRsLiYuwCktZoZO5VaSqnMbEW9qsOdBqzKTOTW1Z2bB93hqaxXWjcFnd5mJoRa6tAPJefZfDGfL3Ie3D2EUGvd7kDbG7TiX5EgEkLYWL1aXen4f4NjE+C53eGmOz+trF2QcYhIQpjN52vTVms88bq43LLgS+LCQXi7heDXRjuGl3t00Wbt5vxixbcbHHTh/89/1tkfN/+Sk7+5K3Jt6ZFgo5sTddDTO6fL7EfrfHySS+HU7XVxFmczJosxxhiSg91glXONMe0fXMm1qJaEJBJYghm527Y3rjBIxrAB4qbJw01Lrq3PIVxr6V1zSxVQrUTsbm7Vq1c319IyppsA3ZZ73U1rbQuyXoqZqlqL6B36taoxsddacq61hCAON3MCmFmCDMsTMwsxNvW8SYpuZuaqWmrZWSxiTEPfD0NfSgkxxhA5RMCtlPVqSWCREGMCITC5KTsnERchMwAi3CJHjCmETUtHtM5zRkIhBGFJKcFBCjAMVt2y1mIe04yYDXAzNVfzBCaS6mQQMBtaejV3O3tmfjLYSul0Xe+e1l98efTzz+7/x4/v3n+87h0GqkTqcBCBx1yIZ/wq+FupPgNg5t39nYMre3t7O3fv3H/48Oj0ZK3qMcaW5cxu5CBikSfm7ASIjFZ3bBJa3FxJW/FZSwwHHOdX5bfnelzf34SdjFFmBnMnA772+4gAoRaPAbgTNe16DPZhEBMxAc1w4M4gB6N1xayV2VIMIcSUJDARTKvCjAhETuwiJBhTy4kRgsBAoTsdcnFU9f/x//qLv//BjVd3RiYmJiYmXimTAD0xMTFx+VAXpxBQipXY7fjOQgd3LR0nzVoG7bqZSMi1jNHJamquaszkjlpLq9hVMziaiXiMs2ztjGKUzNw6JxFqKcMwqBPCUDh1VH9wc/fBcnXcLx2kDj9LbQSAWuvhw8O9A53NFucTM2qtzGN/c1UVZuFQS62liigAM9PWfMlxPrp6I1i3vBA2q80H7Q5vbauAbfTz1gQtxEy0u1jUIZchv7FiyxvJiyvI36Mu8OZLut9Bg37pYR1v+CH6bmwP7CWVpc6d5adibr/uhD31UemCVPeNx2LM36CXE2HzqhnjjgkGKoC6f/5o/fB0uPPF4Rd3Hx4tV7/30Qfv3bw27wLB1VTLEElSjImqSHBQLbXUmpIMJde+d2ciIRrtwrnP5tVJQxAiwCkwO0xNGQx3N1WrOqZUg1rrP/coUmstucgYtVz6vq+lNKsyM4cYGWTupWQiCiH0/XoMRVB185Pj4/b5RLgtt4YQWZgG6ofe3WazWa21lDKG8Zp13QxALWXd96XUUooDMUU41WqquV1kCe0Ki1pLTGmxWLgZi8QUiSkEyTkDrRFiIaYQo4gArqoGJ+Eudu0Ta3tvM+FmEKcQBeIcxMxrVdMqzN3OjgIw39+7UmspZRgDvYktziTMrsyu/ub+o19+/pv/9+cff/zV6ZdH9bTUAnIWa/3vVDEux2yNt5dihL4EYorv3br5zvXrZnb48NGD+49K0VHFZTI4bFxzj+HinN2bw6BZlx0tpyVSIOaxjozG+J1t9plvlOsx9mwTHU5j/gZV9lZZ5qbnD/82t0eIAnEgIsDc1ZXJicRs3AtzqsCmdQiKuRJFiXBnoq5bpBgI0FIN5lqISYS7LoQgwhKjhMAizORm2vdqJO5hlcvg1OXhv/jZ7/6vf/7L13N2JiYmJiZeOpMAPTExMXH5cArJV8quauuSzbmZTUSYE8FZRDbdxltH9ABAtao53Nv8hEASRIIwkTna48zSKsJFJKUEa3PmysQszFGIcGURf/LBzTuP+k/uLel8TuCmt42qHh8fz2bzg70r69Wq74c2lTd35jMDjjAXkVKqmfMIjVbt1lYRIMZWs27/LaU0rdnMW6Qh89bZvbX5jDL01lbGIZgZNiL1xNfjTwVWfuft4NXrg2++Bv1Mnn9wnk4L/V54kw/spdSdN6p5s3mSj6LPxae9yGc7ayn2De91tkE694c39fA94wO5w8YEBli1qnZHa/ns8EFvv7x79KPb1z98/90bV/eu7M46ZifUJprWTGuvpTR/czWtZl1KBDY18gpVzX2pxWFIsa2Jmqq7E8Zkp2HotV23xoZtVEpm5lnXlVJLybXlKcdARLX6MBQzCzGEOKumuZR+3YcYO5Jaq2ptgVREJDzOv7xd8tSNTUDEBAlwr04KAVNKsV310nwBIiVhCRAWDgQQc5BoZjlnMAvQhS6EECS0ZI9i7k7ixAY1MgpxFtsCLbfOEKOv1iW22BNnHsOmVbXknHVwMLNE5jQTJ9HWwlhNhINIjNHVCAgSCeomIrGbLeJ88fB4fferw0/vHf7qy8Nf3zn84sHRo2U5za6AETnMAXOc3Tqc3U1cvAa9TQ7obc4YEUT45s0b+wf7q+Xy6PHx8fFpqUY09rVw8nbXQvD6VBXX+ZsZP7v5aQ7k8cFNXDTo3AFUdQDmRptVfgIAM1WtRWt2rdiEq52HgcgyCzEC4uO3V4thY4y1d04wQBjgdu823vQJsxDHIMxkrmxOMCIEphBYmEOQmIIwmKndh7btcwjZvTiZ+iK+99H+ycs8GRMTExMTr5dJgJ6YmJi4fPyDf/iHf/ov/7tdprXZ6XLVhVb7SCxgZkYgyMYdQwAJMxFKLd4m2MxCLOPkoBUbbySxjcjLzEGCk5mZqYUQQowcowAHO/Gj92/+4vOjLt7ri2871RPGXFFTWy1XJRcRcbXc933fkwi1Wt9NkoYyU62lWIvjiCGICDFtbWJE4LFmlIiolUW3OTwzN7sZQG0ix8zuuslDZGbGZkomEkKIVavpG5t7+rbyGrI4fksN+jVb7b7V3r6ApRV4NTs//Z68Ws6O77cZEc3H6Oein5+wT29N1Zv/XtCgtz+396Q3MRf/qR1q15TtbjtOKk4frj5+sPr5Z19+cHP/7/3eh3/nR7c+un39nb35PEokwF3NrNamW1Z1dQNBori6DlkN0JLX61KruWkOqlpLzSUDLjL27x2Gda1m5q3BmsHzMEgIe7u7pda+71fL5Ww+293dm806EgJVMBNHkWgggypISEiiVSvmVa0ZoqWbtRVUjtHNjNSYSUREYuxAcHNml8TzxdzdJefUzQAYB6YxQAMOIupm81pr9VMWYebE3HVdCEFV1+v1ar0GyF0CBYU7c9d1bm5uSaRd/UvJbckZm+Z1MaWUktZK1NeKtmshxdh1HELOWdXckVIKgZmgVa2qjwvJQhIRZxZ3Pn3w8M9+8Zv/8Mtff3Z/+eCkVMC2g9PdXP3imD3/00tZB31zIXIJPF/M3nnn2mIxO3r86PHx49PVUs2J3KqDyLkJ7+SO4vXpjbQE8VYttsl13jqeLx69bQcOIm3fIQxv4RvkDtOqVWsxzW6GrS69fTkgoCRhFiObk1qrfTM0qRuOc6tqTkwEkaY7t9KDwCLclOW21EFBQoohRuHAIYYYA+BE23s/ZiJKna4GOFXyx3ZyIHsv+1RMTExMTLw+JgF6YmJi4lIyYxpc2Tmr3Xr3nYDdsj6y3JM5d10tWlW7ADU19xQSM5s2j5fWWjgGESmlqOpmWjIak1XrMAwiEmPkc2qAu7d6yRRw7cri1rt7N9/ZqYdrW9cndV1ywEzX/frk5CR13QFz13UkLSfQt3GEzazTdduKcLi7mjXzNRMTj7WkzROdUmqt4dsWhmEA0MKs20dgZgAgpAQAACAASURBVBFr22Uip3FiFmKIKWo/xUC/CG/UnP8FBdZvq0G/Tt/0BQn+xY3hL6g+vwreOFXy7WI7qi8eZyLyVlk/as3bgNcLSpA/oSwTXYy/f3LTXzfm2vfjc5/yfeHnpfGtIukAwYdNv4HHPX715er+o1//6uMvfvze7k9/9P6H77/3/q2b+/NdMaurU4IBNeeeg4iE5eqk5lL6IcC91rxem6Oa5zw05c7NW2Rzms1CDMRhvoghBkIL26VcMossFvNS6mKnHFy52nVd13Utx3m+2JHQtl0Xs9nO3t66X4tIjGneoqUAELNIDHHIWbUu5gt3z6W4OxOFEJqfuuTanNfNOtrNd0opZhq7WWgrtURu7k4hRkjozB1OxCnGEAIzG7FEjWYAZt1sb39/vV7nnLVFLRBLiF3qYoyPjx+XnEHezboQQimFAFUDeDZbzOc7pWYAXdeB4YSd+dzhZqZmZqrAarXKQyEOHJLNuvuPlnc+/tVnXz36i18//PT+8aP1+iRrD1gbrVs/++b8bldEzlZT3t5vIAK19n/M4cqV/R+8/97u7t6Q8507dw4PHw390KXO4OrWWmCMivKo8V6smGAiFtaqDmyWJS60cjy73drWh7mPC1lOm/+amrUKAAOo3apdiOBgoo6l5am7jWp4s2e3mzVhkuZchkGEWURCFBYiqI63fgYKEoMkQRROQUKUEJiZwHDXEAMT3JREgoQU4gDJ5uZOg5zU/Ed/+sev6txMTExMTLx6JgF6YmJi4lLys//yn/7Jv/rHkAxLtVaJUquWPHhRstKCNwzqLSKQnJlTSu5Q1VI4xiQsVc3NRqkDsBY2OXZpopYCqdtHa4VCyRUkCNcOFh/cvv7o9N5yVRXAk4KBma/X66OjRwcH+zGGUgXAVhH2saq5dW7nVjHaVGbyzYSJjMFO0lKhmy/btkGDm1lVq5XeuH98q9S0BowEcvcQQoop52z05hn+Jl4Ov71o8eaobxNvOc/LATpvb96UpDzzic/5q7ONPbX64Q7fREcTbcXA791t+vQHofMPbw6KO2gs7iH0FaXUk9Xpco2Hj0/uHpYP7i4/eP/4w/duvLO7WJDPAsUgTkoEuGrNWivQfMlROpCDzMDMLDEEa1cmMw4BRGbGQSTEEBJAbg5hEIE4djGm6PAQQghhzIwKQszuDqaYIjMbTFhCCu5xvEiBCCwizmQaSQRApFaNxCFIcyKztB2xPGSW0M3nHIJWdVi7aEoIY6kQk7DMeF6rApAYWZiZY2AOkmZdKUWCkFDsEgmZmrsRSEIgISeEGMAURGKKTQGvtZpqi91qZUnuxixVi5oywbya1lyKOUFCNqxdVqv66PTkwdHyi3unX9w/+vLB0ZeH66N1KYTiUJA38fOp07xdAN+uNNAoVT+xPHI5ubB0RLS5CXH3q1euffjhhyHGR48O7937anl6UmuRkEaluf1Lvll52dy9nDuEdq58zbf9oM9Hc5w937ePjPvgDji1yrXW6NIVW5F6+5JzjnR2kLmrmRpM2cYPxWBhicJBqGV7cBPN1ZyJCCGIkAtTCBSFYqDAFIRESBhMYIGTOwwkLCIsLb+6FB3MCthR7z0admbyks7LxMTExMT3wyRAT0xMTFxWXNwlYGUPDh/szFM9Pc3r09oPZbD5fBG7qCghhBiT1krglDoQ3D2UIBLgFKqa6ThJMTOtbW7fdV1Tckspampu1QA3NVOvxX3weGV39tEPbv7q06OHvt5Mgc5r0L5er0GPFotZjFG1jn4p8w0tlpCCSHsvNYN7i55sPRJZRGKotTYROecCIITW/8abd7v1NjSzFje4eXN39yAyCtAinqL0QWt53Sfp8vEaQjO+Ldv9eb4Q8eIa9NeoXa8EeuqPL0tOeQPP1OvkTTDtfut9aIoOnVNXz/KLNoLyBTH4GxPBtwtv/ixBejtKfGM+hRMYNMp8Cm/LjS/+IV429LQZ/LzJe+S8MO+jH3T8dA9XOFqVX925c/A3X9165+Of/fR3/s6Htz+6efXqTtgjnnWRSOGVXIMQhyQ8I4oAmam7ElOXUuqSVgVBWHLNfT8sl0v31kItADAoCZvZUHLXpRDF3YjJydG8p+a1ZiJKs44J7koEYggTmNWs1tpsy2rGIhIll+wOZkkhhhhEpJ3DkASAqQ05Nzk7xGRmrWjJgRCTalVXg4rIrJuVXMxMpMVgcJAgIsx8enpaSsk1t3Bqq5skB3eDaR1iFzvuRAQAEXWpKzn3676Fc5lVEoJxqbWUXEpWzVoHrUOp5iSU5h53egpfHj/+s7/69Z///JM7h3o6eAZAMELxZmgnXDjNz/4upCaKclsUf2alwKXhqXUdAjFvlF+/du3aBx98uB6WR0fHDx48HPre3atVgNzaQXMfR/pTodi++QVw5yAg2qzrX2T74LkbpDFW3QAip/GbYUzGaE8h8jGD+dw6AMG9mlo1LTx6CIiJmDmOAjTDzaAMh7lqUVhMIaUuComMic9BiJvwDYUbwIC07wGHcgizblZyrX0tWZcgdeoDrl2Jh0fTLdzExMTE5WYSoCcmJiYuKy6M7O4Yat3x2bV3b/bHKa/WWpqYXLNmNTUzLR44zbt5LaMQnIdc65hHGaO0aA4QxSAE3orFbVI6tgFsZbMGuDN0f5Fuv7P/zp48fIRHw9NzSTetOQ/DMBCxCNdaah3jPpgIYx60tEaJAJqzpZUPi8hmcsMk3h630TltAItwy+JoMvR23r4RYgBvbja0TI8QQtcl0zJp0N/E9ky+LGnvO+ukT7/qRVIpni9WXFop4xm8dO31Eh2cN0R8/y77MBphz23CnzAqnv36nclJ7nQuhqMJ2Ocr5LcWx2/KrCGgRXY0uWnUoc76kL2JPGP9ibZlO4C5G6AAA48HKw/69fDpr35979Z++tGtgx+/f+2jH928ejBfdDOhCgcTM0UmYWa4MTm3qxBAQk0aZJHUJVCLZWar6oYYA1HXqouYN25eOr+XiYkBmBkB7hbczWwYMril7DatjYwd7sLcpVl7tYg0e2y75o6qo0BEQFAzYWnhG21FVoJULaUUAMzcpY5AVetYuqQKgJiEZDabpZTacDIzEvG21htERFik73t3E5ZSilatJY9pD+6mtZaq2gIaLNeqqgR3RGPRgFWujx6uPr3z2af3jj+/X+4enTw8saXSQFQc5O14bofq14nJFxdZnlx/eGNH5osz/k67u1khopTS9WtXr129GiSeHJ8eHy/VKM5mkpg4NrnZHU7mYxhz0+TPbbHVpWHsmbk1l7cqM3rWQTvLgB4XwFqtmzNQaq5lDORwV5z/jnpK/yZAWIQQRWDGDgbadhgtXQRMFJlnIilKFzkEEqEgIJiZlgpJkUXAIBEWJmaWNuCDVj3uT4ahEidzrnB1m5/slJT/9X/885d8ZiYmJiYmXi+TAD0xMTFxWfn9P/ijf/uv/rHvkJ5YrkNM160b2IgSDXkYCkUGC4PYrDp5m/80vxWxs4BZWNjBjtaZMIQYhbnWqqpQBQUiUjMmMrgRWEMg60iuxFRdfnhj78Hj5dFX/dO7Z2a1lNVqHUKYz+fN/NzeUZgBEHjjxGNuCgCNNsAWftmcNW2+3fINzTzX0mbpMaLp7CKBiMyUWgckIms518QA2J2ZXWRu7eFsX2MUmngrePMDRF/WHn63jbwh0u3fap55Dp5Y9nn6GU9Gu7Y2X9tXPSfU4+tO9rZt2dNv/rpxPJla+0JD2/3sULWnG9yqZ62ny0d37+PThM8f7H9+eHLvJN++sf/u1cXOLM1T7CKngBgoMQtB2JlpFGcJcNeazZ3gXQohCIGyVmdnYhYGoBu7qGOTJTXmSwiHQIBZGdstqAJgZjcn4hASICC2Jru1qIFN1zhiam3biMjU2qUwdQmAuxGFdt1sl3EiEuYUEwgxRhYOMZJwS6BuV0wCtdogYWZQzoOrtgNHreaJQHDTompwzTnXUhxoQ0uY20W81qrqRqygalzMq/lQcf/R8f2j5b2j1cdf3PnNvaMHxxgUFVDmCtImdI75Gv6sIbodwM8YeD6KoPR1T/h2w+V1s5V6n9Rxm/sY1KX4/nvvXb1yYGaPHh0fPT6pCg5JIEDrljHeCPl46J7hgKa2es904QBcEKB9u1ZF23/GJS/abJcAuMF989+Le8/MkVg2vaRbU8HWx1ocLUajmamFiJgjcxLpgsTAQeBQd7gzMcb+iC1Gh8mJDMRNQFfPdVA1rVaUOMaiVYPk6kFyzOklnqGJiYmJie+FSYCemJiYuMwkonU2wrIv69XQ3MBd15GE2M04iLnVWsUztZbiEkggIvOFgKiUOgzDus+AE1MIQkzEFGJo6m+zRcN0nOUIs5EAM4lKIQT96Yfv3H/cf/zV3TZTIWIfqzgdDlM9PTmZz+e3b18jovV6LSG0LklmBmvd1711HWwT75anAYCFY4gxxmEYWhIIswDeD4O5M3OI0cyGvm+maYxNCCWI1Fr7vj9riGOmqhKjupVacr92bQ2QJiXuTea3sU6fl9VeES+o2X2j4+9bvfC7ccFg+B0O7Dc5a18fb86e/FZ83eg5czH7EynPT8hYY5rGxYNwvnjhmdsfu9qdadlvyGG8qKA9yTOESz87DBs3NNAiBcyhQFEsezz4/OQXd5d/+v99/sMbez9+/+pPPrx16/rBtb35ld3F3iIhhSRGblbMgbZ+WcfmhC7CqYtWi45BVWREqq6mRVWYAS81ExOLAOzGbpKSMYub9UPf9NydxXwxn1VVCWE2W5iLOatjFJ0JgVlERMhhqpWZmdjZt/11Sy3uLkxMKKW0a7SbppTm8zlx69ZgEoO4uI3K9Ww2M7OaCwAmZuaSh5yHwNLc1kO/rlp9bL5gptq6FJuaVlW1EKRdWEsuBpI4o24XSEfHq6N1Pjzp//TPfvnx5w8eLT2bFoPamJhRrWU7bIdh6wy8Odfb83puCeHpU+5P/PDdvma/L84+6pOLjb79QLNZ98EPf3Dl4GBYD1/dP3x4eFIqUhSWAPCYiDGmzGzjcXzbIKMh3NRg8lazpsbMbeHh7C3PAWCzzOGtsQfB4CCglqxarJVE+Ln93ZBEZiEmDuJO7mQMuNXaxRDbQg5AbuwUWFIMSSQKB+YgALTk3hgeZTabhRCEiZhbNYI6TD0w3FVLXi5XDoSYqNs1Cj2Zmaeyo5z/+3/37176qZqYmJiYeM1MAvTExMTEJeb3/+CP/s//5b+aI4F4NeQUO9RSVGut1ZS8OZyYRJiYRAhuprkWYg4ixBRiJAky5idbq8omZjdTt6IVgITQopsJlLoORKUawXcj/84Htz9/MPw/f313ABcnNTu3dw73Ukrf96vVqpSqama5ltrm1QSCEzMJS62VhUHk5sTEzFZLLiVkKbVqVTUNIhsftI0h0cwpjaaYVnc8TqTNHDCt4/R3M78W5i4lLdnMcC449bWes0vAW6DLXwofNL6/nXyR9/1eXbHfwJu5V9+aZ56GZ0RwtMfP/fEZsRRPPv5siM5Le28BT36KraBJDqijqmfTvupw9+RwWT65s3znoHt3P964vnf7xrUfvPfu3kwSWx16YY4xMBHUtBQRuDCstGtH8+I63DanINfcOhA6UFW1FpGUYqdqqi5Ci8ViZ2dHS+26NJ/P1NRbe0MKLTGhRTWLkJuaKksAsRPDzMlF2E3NPcYQo8ARRJoqSUwgUlM43DY9egGzUWu2qqo6OMws51xLFaJZ6oZ1n/NQiE2bObu6G2BNsXR3NXMHSzAwyKjrWCKInPJ6KKfH/cOTx/eO1p/cOT1cleNc73x19Oi0rgsbxDfqqj/zzHzH09qSo3/75KU3gE2DDALt7e3euPHujVs3iOj+va+Ojo5Xq76oCzvg7lVt7Am48caP29iWLJwtIRrc3W00Lbv5k/dgLamjRZ+1V5i683jjY7TRm83UzWAXjepbfzQ72B2m40keDdROgDAn4UAkhECIzK0kzd1MyEmCcJwtiF2EUkohCAGqRYuZibsBCJXIFV5TEJYQYufdbF2qQWqpyqu5LV7RmZmYmJiYeJ1MAvTExMTE5aZwfdid/GR56zSvr6UrHDvLpc1jTJVZiJhYQGQEMLtbVRVVZna4BIkizE2arrVWMye0lAp3gJk4CNTcvLmViankAtdA4b13r79/8/H1ve5o8NOiahfqyL1q7fv18cmxGwCs+74J2SIMkBtENuo3c7OESQgiXHKzffG2bWGL43TzOlq1VEJgptbYEOP82bfhoNoSEmksr1Y1uMcQJARVNdPRlPUNAvQUWTDx6ngR6WQagX8beX5MRwt+eNoE/fyx8mQN/5sv2r0Q5z7FWUqtb+Q2c1dFOS1Hp+WzOye7Ha7v0Y3rez987/HvLMvVnbSIxFZ257O93YU0GzMsCow990ZAqxwy96rV3EFgllwzgBhTW/gspbpLCl5Ldgel0HWpS50ljSHEGKgi51JyJnbiCCKSQASGFK3D0DN1xGS1qlaQp5jaNS6kJMxEZLW6mau2fAytdVxYrWbuBFJTABJCKaXWOhCbWam1DAMT1dmsX69KzkxUaqmlNCcswVmIhUnY3QwsEsBkbD1iLVSqHS/L4ePlVw9PPv/q0Wf3Hv36zvJxry11y8AKtjG4WQkYo4gJv40ovHE9n+VDXFLOyfEbAZr52vVrt99/b3d/9+GDw7t3756enuZcDazmIDO3WrWleIOImbahzechoIWJWVONiVgYZhduZ9zdVWnT6rm10RAmIntCgHZ1s6fXc1rydCASgMyJjEDkYBqzQoQQGFE4EITAgDAJgcwAh3PLUU8pEDnIRQJA7qbaunSMN29uLuSBvUspxCihKywrVPU6aI1ifzTZnycmJibeCiYBemJiYuJycxzXN46v9bA8YH9ui8Wehz7WaFqLVic4iBxqVktphhqJwdyGkplJGAS16mpqWgC4e8nqcCKez2cA3CEsbJxzVlUr1ve9OcApdLNrBzsf/ejdX3x2eNqXbc4hME5fTOvQrx8/Prp69brE8PDokEApJido1VxyYGk1pK16l4hFhJmHIbu7CG9pUnItBUTC3OfBzUod/dTM3KqHW/xlCOMFjpnbHMfMyI2IYkxunstA3yg+jx/jbxWT3PmCfOejRE/98fmj8Hs8HV9ntJ34rXgR9/tzDv22Iv9C1MbW2nz+tZtADz/r20dnKa9vKVu3aQvocAMKoThywcmR310tf/1g+ItP7l9dxOv789s3rn30g1sf7MxYc4TOiHLJWQfNOcbYdZ1IAtwMuVQzdcDcJQStZO6qXqtp6bWvBBLmbAFeyxAZVEPMg6xWq5yLqRMLEYMotN64gUspeRjKrGOmsfsCYZa6WmsthUXGvghmGHNC2M1W63XLcGYWM6+1tlBeJikll1rMydEqgyoRDf2qX6211phiFEkhwJ3G+IVihhQjnAykzkqhZ/ry/tHdh8dfPTr58t7hvcPlo2Ndl7ouelKsnI+TwDYTZZMQ8/xIlRfibbgG+dkRIjiDHHAze++9Wx/86IOcy7379z+/c3c9FICIqAUwg0iC0GZl3ZouTE/npPsYQm4OAnhTMvFU2YSbM2y0PasBDh77GfrotHZXBez8tahtkhyBKJEIgQnCLMSBEKjFbnjHHAG22pYcWtCbcCCGMIcgMYUQA3EYJWer7upWpBXmtS8lpsCUgidBDEEkMHN1cyipL2b887uPX+2pmpiYmJh4XUwC9MTExMTl5g/+4F//3//sv6FBfH84WS1Fgi77ThCYhFsPeqIujQoskZlpKYC36QQ3Xww5EYlEwInM1KtWd2MmAGYtrJFSSk6uqjElN4ADUrh+df93f/z+V4f9w6OVMxRkfr5a3EvJx8fHe3v78/liZ7EDd2Y2dxZOlKhlkm76K7UuggBijCAIC1q7mlFHdmLGWIbqIIoxbsINWQKxs6q22ma0Wd1m2mZmcINb13JI8uB4ZmekiYnXzJtZQv42aEBvJi9+sr+xOuNFtrApSPF2OdgU8bu/kcPuJbH93GRwB8zhQDFkx7rX06yHy2EeeX+++uJh/uL++v3fPNyf89VFurY3e+dgZxbjkJcxLcJih0IS9ygFUqqWWmsKIQRxBCKLgZgCO4TGBVNiJofX6sylWB5QS3G3tiILdxC8slZWEVW1WksGEWqt7iBgXbUpg5bzRoV0G6uaGEAppWUEM/O4rGBCzE6tkEnN0NocGjcbaiAWJ1VDiJFjrGpMLBJqvx60nCxzMV/l+vDxg6OVPlrq3cPlg+P1o+X64cnyeJn7DHUYoMRGZw76Np5aMREIb/Wg+s6Ma0MpxZ3dnZvv3bx27dqDh48ePDx8ePgoZxszw5TH57VUjU1wc+siSE8e1nFNwgECMW9T3S/k9oxdCjEK09S6PtMmT9ps/PfpGyHaOKA37S/dHW4EELg5oNtNphCxe2QKIlEkBYlBxoAOgmo1M6Exaby12AS87TXQQtgoRk4BnVAQEYnEsawGrwSS/+GP/+I/+9G7L/2UTExMTEx8L0wC9MTExMSlhwaxxVoKTrzX4j70e50sukCkDoAppsgsbYqhWge3NjeQTb8aJwosTG2WoADZYKWM/QDdXN2ZOcboMCKadQQAzBbl+pW93/vxD3/+yztfCpF7dhR7wltca62np7kfdhY71w6uVK211qGUEIKItCzLsZ86EZOMkYaAsEgIWltPIzSDc4yxzcyJKIiEGLVqa3rU5PJaazNE40kB2t3d1LQCLUJkO1WbhLaJb+TrRJUXGTzf6jmTevO3i/OLDxeMzM955rfCz235LMTj3N++pYzi3YVcAQPgKIq++uPe7p/0X3zV/80n9w/mfPvdndvvHNy+cfWnP55dP9gdtArvdulAx86NJlKhFbXOuiBMtWYmZ4nkEOYgIsTwsUuBuzV/cSm1NTYgIq3qamauqKZkbaEUbqpwN1VidqDv+1YJpKq1VlVjgqoOOTMxMbFTW0A1olbx0+zeTEQkTAB5kNh1qdZCTCnFqm4kZlCORbpVziySeHZU89FyfbpeZ/XHy/WvPvvy83un9w6HkwG9IgMDoMC4cgEa7xlawRK26cZPmW8ntmwCSWbz2e33b717453ZfH50/Onh0ePlck0cWjdmN7PR7X7WMxAAEwMXE+FbrDMxUfMRE7yVRPATHQibZd5Mx+UKYWIiOKxlPrubQfXZXwNNgz4L92j3WQCDjYQpgAKRMAVH4NCF0KUQWmTMmHxWclY3CAV3ODxGEWGRMHYVAYk0ozQnQRQSEeaoRlW9EoW8/s9/+sH/9vPPXt3JmZiYmJh4nUwC9MTExMSl5/f/2z/6N//8v+5D5dP5CS/3YzpdrlfHfZfCWO8bViGklJIDTkiJm2/J4CwhhuDmpuZqQCVCk4ZLqczbaUQZOxppqaruCDEEDlrLXhd/54fv/eDG7mdfyJ3HddO6HSCMGaUOAOv1er7ud3d21msbqkaRNiOX1manpUITaXVmjswsHEKIIY6tBd206vjzmPVMrWyVmdzGnI22se1znmj+zgxTM61ViWg2X+Q8aNXv88xNvOV8h7WNN9MNPfGq8K/5Gd9mKPhz//jEX42eym1G71luMp766ZIPxK1id/7X8CwtwgAGHMjAsWK98sd31p88LPNPHv/JX927tj+7sje7fevdW+++s7+zEABW553szNPezn4ldajELrIzPOdBTRmca845r1arGCWGJizaJpjX4WARJ1TVWqubp9SJCBGVUuCjguzupSqxBAniqGqlZmISlp3dPREhkFUFnIAmUudcQgoiMXbJc1Ev6kohhtjVUjTX7Ahp3sn8eNUve1+fru7eP1oOuZh/ce/+g6PT07UOFX3R4/WwGmpfUAwK2HZFZBwuow22Kc60GaTbOBin88f6FZ7dS0G78Rg97IQrBwc/+9l/sru7++jx46/uP+hLne/tEwnGgi5yoC23w8+Wz7f/32rQ7f5HRuOzm7m5m6kwM8jd1U3N3JyZQ2R32a49EYExdiZUb7qyw/XCb3srGhDhVpxGgIAiS2KOxDMJSTgwzVKMQmzWMqmHIWcYwceO0S1czckJEkREiBACxcjuKkIhhBAkRelSDGQMdYVSOO7XGa7u90/Szbm8vhM2MTExMfGKmQToiYmJibeBGir1UanCWUQ8dKVfCjlVB8yEQoiqMx1zJCWEIBxsTF1mVycHMbtSk3FFpJVumpuqUUdjWiDcAFNz81pK0QryhfB71/duvXNw7/iRw2jbrf2cgrJaLlOMO/MFALibOrl704UdrYFSc84A2IQSbqpPfVNJauRum0SOtqVWhkyjV9tGuXnMzTynSjeXEDO1wmQJwcxMn1V8OjHxEvhtQqKnMTkBvNShcN4HTRcyfJ98R4yrh5ea8x+On/XXo43XAAOqoTecVqWVMvrfPDjZmYWrBzvvPOivHxztzedCINe9Wbi2P79xfW8eeRZpFj0JBYJpTTHN56JmtaAgEEXmODb689Fr2nrpEnEQUFB3xNQJC4hI1d3hCCE4oBRIxEOQ0CXpIJ3DRcJsNnO4m2tVYQosZo5amXIFqnFRVsRCdFrWyzIcr8uwWuWcq6qSrIrdP1qfDHY81AdHJ8sh96r3Dx8/XvZ9RjHUc6LzBY/8uev5xUWTjej8jF55Ew0iOjjYv/3+7Y9+8tHxyelvPv/yzp27p8sVhUBtfJ6tmI/hJttV9vOtldu2mvXcAPInFtq3J2n7oLmptoyUTUZHS9AYn41nfg3QZlNCJExMaH7n2NIxmAOzEAuNrn1zo1ZX504whgMCMLE7fBvlwUwiHCOHyAQOQjEGEWZpMR6uCgeUfJmtgovbYtdOTycBemJiYuLtYRKgJyYmJt4G/sE//Jd//M/+UWQmBTFmi7mUTkS15lqzKbSWUkvOuaqZ087O7nw+B8CipVStGiXszBfFcilK5CIswu5ORkQ0m82Z2d1yLTmXYRhKzrkfsnr2fvDTW9f3P7h98y8/mtM5aAAAIABJREFUPSY9a2VzXts9PT0BcHBwBQ5mXvVrd4QgMSbAhyEzk0jourm5l5JrrQCIqNmxQwitrrmU0sJArM3Y0QIQQYQmkW9f0uZvm1BpNzOCMyAiVbXv+5xzqdVr/V5O2ZvK65QQ3uQIlBdpFPd1r5qY+C48f8w9Zyy+4GD1Z/74Ld/r0vA8I/eosNkmwthBzXLanj2onyzrveXj8OXjODYzBBEOIt7ZS7fe3blxbe/q/mLRcRfQRVnM5wf7B1evdCwcw6KbH4gIC8cgBIdVM/VWlwNnkdR1BCbiECLAbk5EqlpKiTESc1AtpZhbSl3HvHAvpRBz13XDMOScKSLGmGLs+0zV0swfH5+uh+xFJUR1ebA6PT05HfretK7X66PHx0eny8Pj9b3D8mjtJxUKKFCBivHnTc7w1578p//C6VxvPBrDoP27fg224KwW/PUW0Fa9VRWAiNy+/d5PfvLj27dvf/7v//3Pf/nLz7/4oihCNyM3H3OYfcxlPssHA50d31YqRszcYp211jZyaIxFgYJo4zq2cSNe4Bc24knc3VS1RXPYswRogB0CCCEIiXMExyCBOKC1DjFzrPsMMyIXptAEawL4bPmKRtN1a5hIIcQQOQSKEmNgiWNUmplbNS9GErKWXj2DVpoPjlb/8y++fBVnZ2JiYmLie2ESoCcmJibeEoQYpsS+HrBz0C2uHAgVtVK1VnN1GCiEpGqlFAJMtUudO6yUQMywnHsiD4HVrZpBdXQPi6h5MymbAUQxpfD/s/cmv5ZlWZrXt9bae59zX2ONu5t530V49JFKSsoRUg2SIX9ATQChQkipAlRCSMx9wiSFkBCZlEgoQGKYMwYMIQWZhQSVTVRlVUY44RHemHlr5mb2unvP2XutxWCfc19nnbtb8/zZ/rnJzey+e8/dp7Vzvr3W94l0qTOQQjIC0tZODr/47RfXb+zsHIx3HaGaHiwPFouNfmORXeGIKQmzmolZCCFIqLVUEkJMsQ41l1JUa+22men8S4jXT2KGaiJibkZETgQi01pVrVNVtRkTaoNzXVrXJdWy3NdWBH0Ef1Iq6okCu2Nt8k9kAPfnHBwST2xXNh4LD38IPoz0vE4io9m891xD99Kd5z+s3aGAydF4PWPqU70okQMZBDMA7LhdsNorN8v++zfHLt6JgkAUBZt96FNMsQtCfSdbG53Ao/DW5qJPoQvSp5BiCFH6ru/6ruvUq0YIcoeDhIWIHRiH3WlmFA6Qm05CIsEd5ra3vz8MqxCihACSg+W4v1zu7y9XYx6LZnU1z2oHq/FglZdDIfdcdJnHnMuYdTX6YBgnxXlS4X29Ge6/SXGXK8qh8YZP+v03Pra+a9LzAyZQJ9MSImZ0vbz19msvvfTi7dt3Pvv0iy8+/7IUdQ7mtVdrigityzwlOtff5zQLm7I5ZruzqcD5UIeepkxm4w4YHT/fS1E3c1OYwaymYp4gEEWiBE7gABYCO1SVYACc2LjaxdQVJGGuLWxcXzdXQIhjCCJMMCKXYCLKTMTEPCUiTmmIDhgZglrYL2MB5Ww/+H9/ffPV577p3mk0Go3GWaQJ0I1Go3FO+Pv/0T/5Z3/8HxbVwXgYxy4FaIkhpBRHdXMyIjc301KKGciJic3US3ERdcvjGEJkYXa2GgQ4p6zrnJOuanAKIRKLi4HZIQXCfffmvr7z5kt7g965lwCturu3l7puY7Epq9Xa0NnM1I3d1UxNiYiYHOTk6jXNCcGsPt1OI1ENIvUZaH6AORLd46aqrurrAhzUeB4SokKTrwgzBwm1xfX4SJty92h5mO3ZtvkZoe2Ic43fy3X6/O3306tzlxW8V1V4nQpVIswGxwSMhoPBaczwXBVuBgJjESEEOAKjS7LZR4ZFoYubi0UX+xgXXeq7mFLa2lgsFl1M0cy12CS9oXbqCEEOlgfDMJRSiJiISs5mNUyYzT2XcrC/P+YxxOQsChqGcf9gtbN/oO5FPRcdVbOaOY0FQ0a1Fy5E5HWdqAYz+l1X+wFb9KjB84lt53yXl889Dz5riKjv0/MvXHr99VcvXrzw+Weff/7ZF3du76gTgcwMtQa5Wm84TqYN1oWgmpYTqgPLsQTlw71S74Vmo/eqf+OE+gx3KzVRcFafpxU5hhB1QRLXkmcid7jV9jYiEAu5TLJ4dS5nIWYi1MIAMmOCsMQQJRBcmcFCJE5k9SA0dzJTVTdXVqgTwsgYlDP5QOXL77965f3rX2+HNBqNRuNs0wToRqPROD8QfKOLB/vjza+GIQrramszbG1tCHGMKfX9OIzmFkRWqzHnUh8CVE1VVbWUstjY6LqehaNEIipFtZiqei27MVNzIgoUQAoYuasXtxIkvHBh83d/8sNPv1p+9Nmt0y3hRFyK3rmzs7W1vbW17e7L5XIcR+Kpibd2loJIJIiImpo7HGPOZsZ5rM816wWWUmrDKtYZg1UsqIE8buy1SMhrWrxI/SYHrJp1ANC7l1ydMyHmLHD/B/UTP7qXM+1j4pu5beDUp87aYXPCg+Ahh3fW1qLxCJj9Xyc16h7H+rOkHE7c69ynScejo1Ie5kpTJhhqii9BgTGDASa4gwaVPavC9MbtHEDkVA0+QLRIlCJJIFNM5rwEAsxIDblQlRfhkwLOcHPYXLB8qD8SFcBA5K7uo1k1szaHws1rBTg7kbk5EajG0Nk6S1DmuIXq920Ptng58cpsJO7P2hVjXTj+AGh2Brt46eIPf/j9l19+mYl+8/77X335ZRkzdRsOslJQ/JgK7PMxUe0y6g4yNS0An+xdcDjcTknM0xWf7np4u3uVnu+3CiLSxZSIhcAg12Ja4MbELoEIzAgy+X/U3jImVMdzcpbAKUiKgYVEiBkiLEI+Hc6kTlY8W8njoKXUKurYLQ6KZ/aCHIR2n9/+4/cfuJkbjUaj8V2iCdCNRqNxfohBbutgWWIYJRdysp1lGUdzCanrxxJDiEEAdCnGGNydA3FgUzX3jiAhgOHk4Frk4gyAMY5DMXUDSECSi0EVakRwhzurDh3TWy8/99KlxXbESqc4o8qc9+Ql5729vS51G4uNIOFg/6Bm04CpKsIylyTXahpm6ftuXRE0aSeHCTumpgQCE9GUNOVuk0awjuWZ2qshwkGmSHpVJSJVSzEtDw5Wwwp3KTw6wTNW3fV4OZGDdD/H1nt89tu/5+jb7j+ARyiyPOQh9Ki+8ZtUOjaeCo9vD/mhBv2ED78zxf1P7cOfrg14TxVI01Gvjsm/YjKQnkuLAYYTwIbRnHx6vX5NGCAMYrgd/oNDBDeYQ2dJcP0vDR1xyThxlayKM2OSp3FSGZ0dG0BzKPC6+r1Kz4dTEX7k/feAjm0h8lkOP3z1eGX9k79gPgwPOar7f6M/3JC8piWnFF55+aXf+Z3fZZZPP/vs/d/8ZmdvN8QQYnSQmYvwiSLlo2XQU4mzu1u0tdsGExHVLrXjNdBHB1+71w4XVIuhzSwPq2m+YV1HfWQ/Ug0MBJFzNfkwU5iRIxAzMxOYIIzAcFN2D8RREJgDUQycJITAQTgIEYEYIhKCiJC5OVAt3axoGbKWEWYhxO1LW2mxsbdaqZqzbdzc/aNfNffnRqPROG80AbrRaDTOD7/3B3/yv/53/87q7YOrHy9GUzZz1TIsAQ5hGFfj9vZ2SlHdQowhSFEVEmYqSkQUYqymGEdsBWvXpKAQDCzCkkCiubgRrD7dEBE050jyynNbrz239eKF7rOdrG6EWr+zDmYH3A/29mNIL7/8ct/1wsHciZmjlFLMLIRgajWBkIVFRJiJaJKdrZY329xj6qpaa5/nZzZ3d2YJIVTjzpqubqalaAghBKkCtJnWR7gUk6oN4+jQasB438fLpkE/WuiIBnKfbXvi9cdazPuNd/HDf93DTHU8Eq0E7Yg9szzhHfMwFhvnUnU+wr229113xX28fQ9bCmZ/ZtCRBdg8V5r12AQXYc77+5qDfuBl8ZSNwjSiQ8OV4+WuDrK5pvsh9dRTX3zymnzE3OXMqs8PM7CH2R5HJwjusxwKUS5duvDa66+9884Prl+//tFH165dv17Uu74PMbiRmUuIPE+fT588QlWb64vVf4xrDmEVoKcc5tPD8PVOWte2VxtpUy3D/daSiIS5+jubw83ItJbMC7MwTQI0IRBAzu6JkYRjkBA4BYkhhEDMxEdEbZpnOdQ0q7lBs+bVwPAgxMxd34OJJZiWN/7iV3def/5Be6HRaDQa3z2aAN1oNBrnitXl8fKXiV2NaGtjI/FW3v0KDjNb7u+XcWQRh6e+CykZpgh1cyORw0oZYrhZyQSvpTB93wNgChw6gPNYbBx1HKwUdzAxlVHgW1343mtXfvLO6zv/6tpKRxBrzVAC1o87wzjs7+/lPKauSykNwwC3yIkC1GocvJlb7S11d4TAzFNXcn2kdphZtd1IKVV5GlONtasqE7Hw/PiGah7ibjmPpdDaeJqZ4HA1B1iClRoHRbND5nlXY84KZ3A737Wg7OE/8iS5l4z5bQ7g76Jm/TAm42eFWrTYsk/PEg8/5XOXT51Q8+51/sxVxF9vv9/73XcZ88Mv+pvozg/gDF7JHx/8wHeYewjxBz9454033hCJ1z/59MOPPx7HstjY6rqNnIszBWY/lQjKzO7IeawGYhITEaa5dp/u2VB158Mi+sPryTrPcHobkZkdaxur5ffup4/aekgJ0aSJz4X6TCRMwhyEI1EgsDu796lPUaJwiiEFCYGZSWg9IiO4m4/DOMJBXqwUK0WVEYRDjHFzo99c9KnvKHW7w0phZuXzn7714r/+4Fvtn0aj0WicSZoA3Wg0GueKf/AP/vRf/+E/utGvInnfx83F1si2Wi5LHl0158FGV9VhWIUUQwgOuDkHIaERtcRFRKQ+irAwsRALM4cQY0gGVgVR/TFziA4Cc88ixJ74tVde+NHt19778MuD1TiYo3aiEpubwwEyK+O4vLNza2trO4RUSjF3FlEzh4sEVCnZHHA1s5yPOhlWM01irkbOVU52+PS4Y26mtSjNVOvTWn0LT54ctQDaVY15Ut9FJMU01Fz4iWfqWbpxHx5GjT2DR8u3GdJ3Thh9SEuWM7Ne9zBnfSqchTGcMx6yj6NxTpn2c9ely89dfOeddy4/d/nGzZsffXTts0+/yEVlyK7LnAtIWATEd5lIMC+qk8VJ9cFQnRMFDy9lPt1hTSXSR16s7V8AyOkwt7AK0DXz8Jjn2LxIAgQI1dHMHe4EZ0IQisKRKDKnIEkoMUXmvk8pBmFiIgcVcwGckMdRtfa0CQOlZMBADnZmShy72KWYUoh9F/u+C6nbHcfBdXRjxnBh493HsmsajUaj8ZRpAnSj0WicNza8+/tfvfhXV6/FkPqtRd8Fv/klDszITdVKGcchj6swhL7v1bzkkvoOhLGMEoKEUFVgIgohsAQS6bouiBDctZRcyli0GBwsgUWceWNDlGhQe+Wl53dW5aW//tXtnb3xQAUEZogUhbnVft9Shltffemmly6/UEoupdSQQ2Le3IrE4nCQqWkNSFwnDRKIAQkhSDB3U82l1DRCFvZJfcYUl6gGr3U4RkQpdUS0FqDXOfIExBDQeS55CoA6U1rVd55zUEv+gD7rJzeQZ5ETFr1r5fab1auueWon+BwwBhxZmSfDaYsEP/WGdjQ3Gt8aB7C1tfHyy1ffevvNFLv3f/vBxx9fv3Hjljv28wF8CQdJ4BiZwwkPaJtNxioll9oZxkzETHOzF6qx84kvPswzdNS7JqJ1F5o7JrtxHDnbj9zvMCCAgNgBN3JneGBE4SQciKJwF0KfJAoH4thFEa5y+WjmrtU27WB3bxxHM18suhgDuRIZC1KKXYpdShv9ootJarC0cPZyUMahkOdyl7VqNBqNxnmhCdCNRqNx3nhzeelfb+wW6/a1hIPVxQtbWxcvdTGUYeVmpZTVakD1miDEwKnv3L1o0VpvnHPVYIk5SKzOgzF1woEAkRhDSqnvQmQWNScRDnHUYqYJ/sKFzXdef/nv/eyHy5F23v+kwNWtulv47Ehp6sMwDOOopkRk7svlsqgCGPIIh7mZu8HN6sOSEybfQyLyYXCHEAEwc2IwM8BqamoSJEoAghVl5pS6WonDLCLMtXTapwpod7eiIQQWGYbBVI8UQT+zPNDdsrHm7G+lczmV8u03+9OZZKLJWv/Idz/0QB7hiM/lMdFoPBHuevE5dkpVzffll1/+yU9+0nf9J59+9jd//Ytbt+8QCUuYEv5q+gWLsNBJF46wdnwGQVjcvZTCzCzMgPlxAfouI3LA6w1Tvecxs5rw4ep2cryHMFFgJgfBBRBCZI6BI3NgSSFEERF2p5K9+DjmDHI39Sk+xAKRMENdOHRd7LvUpcACZg+B+kVaLLqNvtNcyE2YwcRdPw4DhFHUWeH0P/7fv/z6+6XRaDQa3wGaAN1oNBrnDXr33T//w/8837gSX/p0P+VtSL+53YlY6sytlBLTUGPPx5LXzydsxjGZmprWkmR3KmpaNOdcFEwZZoFDlFDSEGMnIY5FHSDmrNngEjhs2IbQ2y8//9sPPn8Pn2hN1KGpL5TmOMKSy3K53N3dFQ4pptU4VHnFrfaJThU7wuxuAEntPJ1qlokYUhNuyJiIiGt0O4h4Dmo3EDOHINUGmmYmR2kQMcG9fpCI+r5388FW9/VmbdLN16Jtrsaj4jvfl0DrX7NgtJ7q+W6vWKPxrEBHyoYrJ820mSkEWSwWr7/++ttvvr1cra5f/+SDDz4aVmOMHXMA83QnRAQiIT5W8ktEoGoiVm9FhLn2cjFz9WauBdI8Zy9Plsu10tmrI0edtq+fIjVA3Rw0O3Hgbjc5BAhxIAnEkTgyBaIgHIMIMTMTB3OM2Qqc3OEGqMMAm8w6quWaeAoxxdSl1MUQo4TIIpBAKUoXYhdC1gJDYHIRZwymBs+EhSyWunwsu67RaDQaZ4AmQDcajcY5JB9sphe+yKIYyt5yuLx9IUnkbqGmWUvoR2J2YDWsshYz66rvRghjzjmPwzhqKaqmau6ZFEGiiLDBxnFY7u0MN1mihLQac85jzpkFMYV+kSgtVh6f6+X5jbQBDEAhEiIF4E7zU4859vf2h6G89trri42F7wMgZpYYAJibmoEgxFYKHCKiqqoKIMbYdZ1rrXg2mwwOjSVA5k3gtSwa4ziuHRJrgfc6wwdG1WbEzZh5c3PT3ccyQE88na1bVZtM9LU43d9/lLNfO/xd4V5b8rS8edqD4ezwkD7Oj4qndC5T7TypyXVeyxfrH9rFpdE42xxVn0/b2DgAZjKzlBavvfbqW2+/feWll//2b//lRx9fu3Nnp+s3+0UiYgfXC8DU2+VHXXmwTg4UrzPlk6tGF9Y3N2CAQBLE3etNUZWni6q5V1sLqg1k041PNTQrpsVV4XbXdWOQEAXmxNKJpCCCGgvCBAKxEZexlNUIN2GEII4CGAtXJxGpHh1RNrrUp9SFSAQRSoFFiAVUTIchuzJcRETEU9obxlX2wfw1PLfDyz/+P//mEe+3RqPRaJwZmgDdaDQa55Dff/fdP/+n/8EB22bW3d39jbhwy5RXIHJCihHMYA4xFi1FixYFQMyLxWKxWJScV8vVOOYQYpVxc85mSoYskonciZiJOQozYgwBUAkUhYZxVcq4kRZXL/Wvv7htd5a3hpIddFxfIYebacnjMMSYuq5TVYBCCGrqxavhhjBHCUzERKrm7iEEZgJQzJkRQsiq5sYcMTseTt9wt6eswyx4NzevAnQNJWSiGEOKacTgWkXoUxaJd/lr4/6cQa3zGeE+B+oZMft9WmM4E+cvgWq3Bx5uQE9+0O1K12g8iGPO8mYGYGtr66c//enly8/furXz3nu/uX79c3Uqqk6lRg46AJqmucn52HWQaIoe9HUr2KGb8/rriMAqgKsapr4KKmYOI2IiJ/dqeUbwGqZhObsZzE7PSBIgRIlDYgksBHaHFnP3MjmnOTmYQAY2BCIndrcYowiJIPBUMZ2EuyB9F/sYU5T6WS0ZTm5MZExSmALBzUfzYnRnuVoVeLavsPtc2H4cO6nRaDQaZ4QmQDcajcb5JLNt7hNHXQ3Drdu3egYNuyIiIUgMtaYlBhFhKTzoSlU1Z+m6IBJAUGNQSinGFEI4WB7kMQMQYuZAMk5PLsRmBqJcBkDd3dQI2N5Ir710+Qffe+n2e5/sDGWsDzBHhlfTAN1stVp1/WJze2sYhqKFiZyIiSE0pQ6SCBMTM5kDKcbqh2hmcCeaRJwqlB8VoGvSYP069+OBPNWwUJXqs1r1RnQDQYKwcl34k9tbjcZj4T5zJ2dEg37yPOXzmjBZt04mrne70LSGi0bjO8LJUujFYvHClSvff+cHMaSPP7r+4QfXbt645U5FVR1EXO+EfC0lz/XUxybpj+jP9e6lOowddYtmVoe7HX7MaooyEZHTpD6DCKZqqlPtszvAp9dBwIkliDAxHKaeYWwGNzcHjNyZPFEQiSlwEGahPoYUhWcBWpgicxSJUSQyB6rtbFqKO4nUlYAUMpgTq+FgubfvVLzYcmFB3/3zP3t0u6bRaDQaZ44mQDcajcb55Pf/4f/8N//lvxdu7N26fGF/ZzdBw7gbQwy1yrfrUpdS6lgY7mTmOR+MQ17FIEFE4B6ZyjDomCUIAUHYDHGxwd0GjdlUzZRiVi2laNFxzAVZQ9dtbmxuXbiIuKFx473P9j66uW/zs1BlLYO528Fyubm1fenSpd3d3f39fTVjlr6PBlebls1EVXd2R03mcdMhj+4uqsM4mFltRK2PamaTxHzCzXny6qjPdLN5IgFmDndmKqWY2+SLPdUPnabpQl+LZ1boPJucqX1x2tzmCQzv6au7x6biiPDQRdCNRuPp4fMla/3r0AC6KsPueOmVF7//w++9+PKLv3n/w1/84l/e+PL2MBSHaQHYiGhOwzhp6LEWoHk9U35EiPbZmmM9mnrPg2kEfuS3WkTt0xw+zNRM7XCwRzRzmtRnEmLhsPaVzmquJnCpWRpEgRCJ+hg3UupjCEJMiIFCYGaISGAWIZ5WhqyWJLiaF/USnAkgRzGgZNXiHEbS0SmDRs4QxLJ4XLuu0Wg0GmeDJkA3Go3GuSXsrfY2O1GQoAtd37OruelqtVIteRz2sFcfatgxKbZqyrlWE88Vw+ymIsIsLEyxcwqSipnCzd1NtZS8yBvFCsjMQcRMdunCxvffeuWt1658env3+q29088+9blrHIbVajkMwziO4zgWU5EQQljl0UwJqA9OeRxVzdyY2N1rojsAZjFTd1+thiOrfti8imOvms/9pOunRqmOiTXtRyRhSuip/olNFnqytKb/Z40TBdrPEJN8dbdOi6d4DvgxearRaNyLY+dH1XpF5I0333jzjTcOlqvrn3720UefrFYZ1fR5Uqh9EoprGbIfW1w99Qzg+eJw9E7mqPqMI31dmLOdiZmJzCb7MGIiAHqoXPvJ6bfpvowAgrEbbBoiAcwSiAJTEAqMyOhZuiBdlCgkRAyLwlGYZbKKFuapucwKVMzJTWFGRE5k5mpGWrKQAyGGXCwTD077N1Na6P/0l3/5CHdPo9FoNM4gTYBuNBqNc8vP3/3Tf/Zf/bvATt9fWKT+4ubzZVgOywM92CtFS9bVOKgq3FOIQURCYDUlJiJzg3vXJSI2pyDOwUlCJOIgkQgeiCAiDjdVdwWBAh/s7y+XK5hu9vGVxcUffu+VT766c+P2fnbXu9gBUMl5eXBw586dcRzHPA7jKCGIyP5yCXhK0Yu7e3ZXVTUTlurgzCBiYlJiJkBtHcUzVQox8VponoN9BLP87FNkEEcJwOGjnpmBVw4vJR/RQ5sw+mi5j9TYNvWzyRNWn5/+YXZiduvpD2jGz9JgGo2zh9/1/Ehd3NhcvPHmG1evvvT5F19cu/bJlze+cicO0UmJidbibs38q01Y4HXtc/2dmZnJHcfU53pjc+Q6aWagWVl2dxiLEBNUyZ0IEgTmaiA3AL4u0j70fjbyGmkIdifTml4Id6EQowSSwBxjFaCpDyEymGrhtBOcmbg6pDETExE7rKg6rHazwQrBRQgGhakWh7NCYickuWQVKiOFDR0PmijRaDQa5592rW80Go3zzcDdpnJYuV3u+41+s+v2+25RrIwl2wGNq6GM4zDmERmEVI05us5GHYZh7+CAwMIBBHOoadrYjKlzsIiEKCGEFFNKqRRVVbgRqEupiz1CTxZ+96c/vLkz/vK9j5aK0VHWDz71KccNwGpYfvHl55tbW6lLYxmLZrUCKLOIsIiwk6t6dICoVmf7uhkWAJhIQiCAmEMItaudmB2uRetSmJlpDviZu1bNTIuCZoNFwB39arl7ZycvV1MX6/EqxSPlgU2iuQ/32Tj3khrp+B/utYRHq1TeXUo49Y0P86UPuSictuC8x6Ie1cBOL/zs1BqfnZE8Efzo9YemkkRfv3JW8LN1kJwnvtk52/j2PKrrc70vsOqdUwXlOmd/YfvCj37yw5deeknd/u5X7336+ecGCykFSSIM8ur3LEGIaspfUVXhWA036sIdEBERqVnJcwqhe027qKMkAlBKOVIEPWVDw2HmzCQs5qZa4CimtV1tvuB4HYwATGBQAiKBXIUoEBgUBElq+TPHwCIkDHcrBiM4A8wcugy34swupqzMDDNT81IyM4cQTYu7cpWqiQiIkbuYwsamgUxIgSHtfvJl/otff/6tdm+j0Wg0vgs0AbrRaDTOM//mf/anf/Ff/2NJB0phmW0jJXAMMblSYNoUXiwWVtTUihYt6oZSlKgMY14NgxYlliAOgpnlUrK5hJWqERGLhFo6LYwaF8gCImZWz6bs5K+8cPn7r734+tVL12/tjwfjqQE6iErOezt3UophczOEUFQd3nVdjDGl1ElikKkx8xRhs07mmb1TCWARJmJmFqG54FlVx3EkovpEN/e/1tieaQFqRgSvwfGzJyOzhJiKFq+R8VS0gYnRAAAgAElEQVQzFM+URnTOOC3KPH2v3plHKMY9/KLOwoo/AZ5FodMfeobhqfIs7prGs81DHvOH3jnVAYPIY4wvXHnh57/z85i6z7748sMPP76zc4eFRYiFWeTQ74KEmd3MptsNn9OTqU6Qzx5oAB32cLGQz9nIxNUcjWcjsuoaPUUPEoyZRQQG12muvw4ZhGO2GwQBBVBkSsQRFEBCJE6BJTAxObm6mho5g+DkTnAL4i4GZzd2ZxAzZstpR9WouarqzgwJMYrEIDEEJrBw3y32Vksgasaf/vNrP33twiPek41Go9E4kzQButFoNM45VsJ4/bULr97cPziAgUshLerOIhtbm12MQaSMeRjG1XK1u7M7rFaqq2EchjETkTiqrTMxmNlNh6EsD5YlF3MLkoqWYVguFotFv0gp9YtFSulA9yAd91tbW8+/cuXij7738t57n9w6GKfeU8D88BnIzMblchyGbrHo+37MuahubW2mlGKMXegCsamFEEIIZmZmbuZHypKrdYaIVAtCYmZmVa1vUdXpM2qlFLibm1bTazPVAmDKECICkHMuZqnvfVhZzvULHk4sOmVz/ezyQCPZh9xKTfd/5Jy14/Oo5cNZG9ujZ5K47mZS32g0vgv4Wn6uYjGTLzb7l1558Sc/++kHH157//0PPvvs8+VyDCEwMbzalLm5m7uoM5G7lpKLGrMyCVUjCyJi0lJsnZjs7u4sHFNY39JUxXkds2w2JScTqNpBmxu0fp+52jrzAsd7uQhgIBB1IXYiYiQAAwyqlhpuXlSLmbsTI8VoVlxL3yUV4gw2Yzc+vJtzYQpRQhQ4q1oIoUtpc2Oz71Kf4qLvx5yX4yhgEnHFSPi33nnrf//1B094FzYajUbjqdAE6Eaj0TjnlN0LF567Q+zLUjZQNi9slJWN42jmpSiBzNzcwRJTv7XNG5tbIrJarYbVQERqrqqmZm4pckwRxFHiOAzjOJaiBE8hwn21XO7v7YkIEZecQ+rj5jb1O7Yaf/DWqx9+fvvTG7dXCjta/ecAERiALFdDXK2uXr06DMPe/r6bj+M4LFcl5cDiavXtOWc3O1EBXUMJa4m0zU2pa53aprIjVqs+IZOV4tzyajVucV1FtPbxKKVWhetDS6DnXz57aO5TSnbiR63QsnE0FOs8Hwxz68WpF9tMS6Px3YDWJ2v1VAacQ/jhj3741tvfK1mvX/v0ww8+Hsdi5tlK9jK9jSYPDi0F86y5myk5kcJB8HpXQsw+JUNXH2hjYYOZmteSZ2Finvw35rRoM4PBDaqFAGZycytFSzYzh61zTzENBewkzEli4MCQ6ili7gYyg1qNY4abw5UJ7i4Ag8pYWDhGEfdACMIhiAQRpq5LXZ+IQUwObG4stjYWm/1GDMJErsZBKMa95TAYZ8+6jxc2N5/azmw0Go3Gk6UJ0I1Go3HO+f133/3bf/KfdPt0e9tHHZwXHEMETM0BNXdXdyeikFIIsRb1xNR3/UiAmmnRUmodTBEJRCTMIUiMsWhxdwK5u6rmcfRa7KNaxpW622qEhauXN1+40F9YxHxQphCeOVmnisEOH4dhXK6EWZjhnnM2s5JzGUuUwKAycyjT+KTn1NqiWsI8h8y7A3Wotf6nPqGZmXttmgVostyYuld9XQMNB4ipPuaZ6pPcX+cCP/WHR8V5VicfA99FSfPcatDrFTtd+3w+V7jROJ8QEc/e7R5TuPTcpXfe+f6Vq1du3Lhx/dr1zz//omR1c3N3NbgBTiLVO8PqTcvspwGaW0CmOXVnCcSTWZi7TZPtGW5W7cPMmHi6ZtS7lmo75pMArUxggpm5qquezquo6jODBCIUCAInm3IPDQA5cdWp3QlgEJEzIEyBJRC6IIsYEocoiIFjDCGFIJL61PWJhUAw+KLrFl236BOD3Ly4hdANOqzIRoMVu1iWd9AE6Eaj0XhWaAJ0o9FonH+6TPu9R46jl93VQS8hdZ0Q55xVtajCTCTEGJkFgKrGvg8pwby6J6vqmIfl8qCUoqrsoQ9hY5NijMJS1eGayW5FteRS8nK5OlgOKx2p5Kj8/Ha6enljZ7Vr5g7orEETMQA31XEclsv93b2iJedRV6aqblaGHEPsUzcMwzAMAKrDRl21w4x4ovpQV/9gZrVNlbn6JHp1gibi6YFu+nz9X5WwazW0rWPlARIW43UR9NlxJX4c3MsD4YFmGnddzl3fX185EfH0QPuFps59M77TB+pdD4n1Gn37Q+LpbJy7fusD7c+/8XXn6566jUbjgazvK9zVyS9c2n777dffevuNlNLf/u3fXb9+fefODki83lG4zp+aypbrjDl8mhkHDsuYq4VGfSfcwYDXfy5dS8G668vt8Baqfp5obuwiN3MirwK0G7zMBmMn0pRJiIWYSUwtu5OZmVbJm1HlaQrMUUSYo6BPEpgj06KLixQWISySpCiBWSKHwCwigSVK6iMJqZvmPI4Du7nDzIkD2HZWw+A0mn/v//nlrVdf+B+uf/ikdl2j0Wg0njJNgG40Go3zzw/+8X/zV//0P7bVPndxb7nauHw5hMCmwlClrPW5h8GTMkvCgLqDAhm5Q0koSicpailaitrUCjq5BJbiXOPVAWFGXATpUtrednUaIAcu1G2kjYs37/zixt5qXIfxzI9EBKr2Gjdv3Nja3r64ffHOzh04QkpQwFHdD9eaMjHXCPgatkNERbX6MjITnBggJhDUDAQmFhEzY0AiEzGIzBTVTpEZRLViqNopAoC7xjTGcX/PSoFPddDn1bf1Pqv17df4tOUA3a3Q9ejbmuj8zTg3h+fpA+ARrtpR1+nHxwmfmZMvnXw30Ymry4k331+Mv+tf1+fYaSW6OX40Gt+YGq9HBGK8+OKVn/38ZzGmL7688d57v75zZxfENRWZQHADUPXnee6c4G6mU+uVzVYa82k6RyFPXh/uIALJoe3YpFY7fDb1qdBk4+FmZlqgBtN1lOE02z6bnxmgsALLrlAlszoyIQrMERSJInEKnGIQQRTqEgfmwNQn6QJ3gVPgIMREpjpakSCgwEI5Fy+uXlydnGCkak4SFmk4GJeOoVB2/eJHb179VVOfG41G4xmiCdCNRqPxTGAlE7NkylaGcRSONA7iamZwYw4gN7cpVJ2YyIl9aut0F2FhSZJMdcr0mx2WcykwJQixuXt9xgrwWg0DYuUwUOi3Lxekf/F3v11lvbnMWFf+rFPegVLKndt3Fv1i8/Ll1WpVSokxWtZqWighsIhUvbiWPJuxSAiBCCg1kwciDKCaigAws/rcJyJa1GEpRgnCLKrFHSLCwjVyR9W0lEmAhpu5iOQ8unsxe5D4fG6tAx4DD9xWbWN+A5qi+DA8ta10lwN6VosnyWk9ITfPgd1nrKfl6aPnzL30ZTquSrcjptH4uqxPUglhc7t/9bVXvve9t3d2Dq5f++Tjj6+tBpXqiHykVavCRCxy9M6kRlPYiRPdnapgXfNK4WBioXVuKdUfziNxVzNTc3KQA0DJxRRwhdvpDorp4gJXcHFjKzBl90AcmQNxz9wzLZgScxROSUQQhNa/kiCIC1mVvB1eTM1VzLxq4GU0N3UlEDuNXgzMMY7F90ddqg8+stju8xf/28e0kxqNRqNxJmkCdKPRaDwT/N4f/Mlf/ck/yj6a0qdffLEhPVa3fVyxcEhJQkqpS11frZEVHmLsY6gyLrFMkTnFVHXKLOQpCiemtLHYcHdzU1VXd1UdBy15XA2qpqDCMcTNq5cXf++nbyzNv/rgyzoqPvLY5QQ3NyvjMORh3FpsjHkcxlFEREIIAQAR1XjAwwh49zqk1HUgJpqk59nW2WvpdH1OCyJwiymFEIKEqWiIwCLMbG6llDIVIrmZEXmKcbFYuJqWMtcbfQPOvpx614LTbzbm+2QPft3Xz/hGO1OcJy3x8a3LU9lKx/ve6eRR7fD19Wrqwa9i9L3qwOcqSMxC2CRLrV9H1bBOdt0fHcN9xe1Go3EvnMirp8Visfjxj3/41ltvdd3i42vvffjBR6vlAA4xBuFAp0/1wyAKiLCauRetfz+CiDChFJ1Mn5mIUBvU6jvXecnTgNzczdxrxLObaVHTPOdt2LxgoylCcQ5RrCK2qRCEJTJ3EjuRnrAhvBkkEiIjBGYGkZMrGQCoA8bGZNZJIBZykJMQS866Gge14gQWca3pIYgb213ayvvDAM0li+yYd//L//Wrx7ijGo1Go3H2aAJ0o9FoPCuY6+Yq7ob9VSmqywV7PtiHK0kkFpEYQ5AqxZpV2ZeIq/rLRA6ogYOwyNxTCoCFpXabMktgQQTUCnMpolnMzYmcYxF58dLi3/jp29du7r7/yZfLAjUcExmnbEI72N+7fSu8cOVKiCHnklKKMYUQ4A4iEXF3NWPhWrPttZgHTjB3qCpqiypz7VL1uUW1Wi5WSbrk4nMjbXX2sKlx1byG/ZgysZsJi4RqhO2Hnax34X7t9Y9sLz5RHrcE3CSwR8UztSW//TH5ZM7Hu50+1e2ICKC16jTFiM1SsvskMPncfn+0gpHmxa5158OC6WNfROufzbo2MP/hXtp0o9F4IPU2YLFIV6489+Of/Pjy5cs3btz84IOPP/3sC3OCwaGmBqLTVwAisuonJoI60X3qPFQzBmwWphkCgh+ZSp/U58PP2XyHAzhczU2PhBweDnoaQ43EIEThQBJBSSSyJOZOQhJJQCIIgcnX3RhEYGImYqoXKCbiYlD1wFw74saSzbRoNld3O8xaJNneupTVB7WVleWSLw2UXxge+a5pNBqNxhmnCdCNRqPxrPB7f/An1/7wP/3xrbf+bOtX5i4MYx9XY1kNbjB1U+26KMKqk1YrEkOIMcYggYSduN9YhK7T6WnG4SQSYkrCzCzCgZk5MIOCiKVEBGJmCUMxliDvvPmvfnP9r38Vy24x91l0JoevdeiD/T3VcvXq1RhTqMXPIQQRNXN3AtRszCMwWTavAeDu1RsaAFVvjXURkk0PYLmUmlK4fpzDofkiAZiUaLfAUmuqmUVEzNTpGxdBf1c40Zf/CDXo1vH/mHhGtuojPA6fGCdPHwLx3D4/K8pz/fIsDftc4Wizj9AUi3pkgfVVm5eJ0wL0kREcXUL9IHAoSE2VkHNz/zNzODUad+Vhrg8O+IWL26+9/sr3v//9XMovf/Xrjz66dvPm7RA6NbOSzRTEoGMWHAQQcfUuY9F5CvwemBMRhOAMdzshQAM1xAIgTJXPPnmamcJ8bfcMIrjh+K2LEJJwCiGRBHAfQycSwYk5Mguc3dzUCDoFRRM5kUidrZ9MqYmHkt1KolDUSs5asmkxV2I31TyMTODAqe8hshyWI2gc7Wd/+YsvXn75v//bT7/2zmk0Go3Gd5wmQDcajcYzxKsHl/4m/n+wYu6rjI1+kwysIIfmMuhKc4FKjEmYQWQKy2XIJVfnZZZhGCDsTMRMzAyWEFLqqAa3swA14KZqIz71eAISU4r9c5uLd15/9ec/uPnXv/z45s6BrYXsGQI5XFVv3brV9T2AO3d21CzOFhwxBIPnUlT1aDIh5mc5ZiZih5dSUCZLaDiqQj0XAx0arXptXnXD5DfC9emOAFXVueQ5hFBKORLu9ezwmOqg14JXo3EvHrkeejqN73HjJ//q1dN+PePmR4sTq8J0eMq5+5Gr1uHZMk3crWVjmj8KOpllWIump/fXHx+pnp7HcGK0TYhuPHPMBhWH+N3+nXJiBOG33n7zZz//OTF/8ulnv/zVezt7Bw5xrH2Y62l1/DwDYOoEEKwUEOG4SfThUIgoTIOxUuDutO7iOpSW61sBprWRfC06hk3OG6cueHWhgThJ6EPsJSZmNqNiRA4zq3nM5EoAMwlDAgkTswFa3T7MzAZzG/JYTInI1OAWAwcREWFH4NBtdUTgwNJ1JDwOZTRXtw/eeeutX3/wTXZRo9FoNL7jNAG60Wg0niHo3Xf/j//i38bBgWy9aEC3daHrNvOYyUxL6breVGvBb5Vl1arrBDlqAyaNw5hN1Y2IicnUqwBdnZeFhWui3/zcI2GyKpRYKJpGeunyxZ9+780PP/5yf/9gMJTDKuSqPoMAM9u5c2dLbWNzM2ctqsuDAxAxcxZxQG3KQnT3+o3r1C6pna0ONXXAbDJX9bng+nBrzC6KtR56CuY61HRgs3tH9Z5OKeUxl5KfPXnmUWnQp7fbY3X5eMh99AgH8DCLelTvqTw7x+EjPFSe2karNq1TbtdaS6qVznOgWFWXrCrKDgA2OT+7H3F4Jrgd9X6u76bJ/BlHrqq+fgtmF45j/fj32hyP9sR8yMLSJ7yoRuMEaw3ajgjQOHrU9X33wguX33jj9atXr3516/ZHH1279vH11XJ0h6m5m9tcjwwQT8bv0ylI84LqLL4IqjEPTQIzYfLMCUHqn10NcGKarg1zKfORexqvk0z1pm2+hBxeMKtQXT9HoEiUOHQcE4UAYnNWsLvUERGYGOSK6v/DowPZ4Oq110xrAHX9MgOM3BkuTAIKwjHGIBICh8DuTiGEjUUZi8LVDEvsb2y8+3h3YqPRaDTOKE2AbjQajWeMfBC2r2QmhsTFYuv5l8pqaXl0VbjlsQzDsFwul6vlmLObMUuMgURCjCGm8WB/WK3GYayS7nK5IubU96oKeAixS12XuhiSu5tq6mKMIYSwGsbiB5kPLvSbP37jtb/c/BdfBahCFeZggA+LmOFme7s7McTnn3u+6xbL1ermjRvVNwOAuWstZ6ZD3ZnmeJ9SyrSmRKC5FBuT2Oyz7oM5+IuZ5+wuXkeB1QVydZWuVdUizEIg1XLvttlzUNV7n1W713p9rarSJ7ZxTlaf3YO72HR+U56KYPcNtvl3SJs7PV1xL9Y+yfffbk953X2a1jo2kqoLHx23Hi+LPmmKc+IlPyI3O06u44keEwB+mEp274E+8oP5IRfYNOjG04WO/4u2DrwQACAnou3trR/95Eevvv6axPTbD/7ut7/58KsbX4E6QIoWuE2fYoCIhKeuLJ/cnt3c4UyxZkvUuw5hWXd0FVV37/uu3t+YGRzCvJ6icnPzWh1QJ6qsnrFlHNUNbpPUjFo5QOTTvQ9V8w0KPcdOUgCQtWRNxCIswpFDDBwCq+lYRiLJTqtR8zjmcdRczA1VPCcWRt/FFFNkdIE64SAkIUrqUkrMgJdclGIk4qyqRqbuyWW8e913o9FoNM49TYBuNBqNZ4vff/fP/uKP/v3t2I3DcncoaZND13d9z26uVnJeFN2+oNVumRxqpkUBqFlR3SCKqYND1VRLLoWYY4zDmFWNicxsGPNytVI1VzMvBLBIKUVBiAvrLthAr165eGPv4PbnO2sPDj0qoQAOrIbljZtfPv/Clc3NjeVys4rFWgqYWY5bKx5LhJ/8nSUEmvpbJ12YcFh+RLTO/aqfqvWEDjgx17dN5hzudSlaykGMxDQMQyn5ZKM78B2Xnh/IY61WbjS+DQ+srH/6cqTfo9z4Xq8/1pE0Go2HpkrGLEFSF65cvfKjH/0odd2nn3322w8+vL27129fcARAakYfVRt3ZhDVhOR6ktf/psJloppRMU1yEzvczEAQ5voKM7n54Y98qnqu3Q7VJw0+VyT7ZI4xT0z6bBYNAAQwIKAAThKFmLTO4kNiiBICMYCsmrXQADVVyxjG+U5I65JDDCEGJgrCKUgMnISqAJ2EgpCEJDGGKEE4SnIW7jZ2V8NqOZjrKKqy+N/+5hdPbU82Go1G46nSBOhGo9F45uhiZzkn9aH43sHq0vYWvJi6uoMlpJBqoKAI4KVozkVVSy5jHiVGdxcWs+qCocQcJIxjLmpwjHkcxmEYBjaFeR7dTN29qKoZE3MYNkP3zpsv3tgffvP5zpyoNZUA0rrZ3H0Yhtu3b124cHFza/vC9nb9Qc6ZmDgc+/eLpkx2rD+rZixyaLRa3wbw2pQaTlNA0JT0ZWpT9uD8QZ9y3Kv7ohMopZJzyjkT0X3Sg84vj1yDbop245GznsM6c0fX/VsnGo3G0+bEuUjr/xNDhF+8euXNN9548aUXb35164MPP/r08y/2V0PsFk4MCIGYaoEwMQGAqpmZV9cyIpodommaEp+tN2BuZmrT900dXe5mk03PDNzNHUQCoekmxdystobBbO09ffz2BwwEokASqklateogImYjUqD4bK+hBhjIPCvgTCQMFgrMKcXUxSgchGPgKJyEwqEALTGlkDoRicIxCCQqx52DAyeo2e7FV9Kw+3h3YKPRaDTOME2AbjQajWeO3/uDP/nnf/QPsbGRR98bDra2+uXB/rC7OyyHLnVdTDFGYja4qhIxs5SiALp+gVkwFmZiLlqISCTUlnEiMphqGceBCEJcxtHMiHh/b3fMI4Xooc+Utp67fOMg/+WvPigZarR+VJpcSoFq8VxK2dvd7bv++cvPLYfVarUSEXWzU+ovM7ubzY4bwjzmXIuGgKmtljA9/K3dPCbfVDp80aymGuKwMnqKKTQAWorBQCesD+76yHo+eJjSzG+mnp2nrdQ4O9znxGw0Go0HcsL3mQg1dJmI7cc//tFPf/YTIrp2/dov33tvb3+pBvA0t23uqlpNMARO8HJcgD4SP4q12Vf9opKzzlHJRFRKrj5mmOfOHYBNk+I+zaY7qGrWBIerzY1c1Wl+uvGppvNT9iAL3EHmRGB2UFYdcp4MqOsKu0ehTpJrZlgQTlFSkhgkCFLgvo9BwLAuSQoSmWPgFCVI6Pu+39gQZiFi8lHpzsE4WClw07J5+8v9S1eezF5sNBqNxhmkCdCNRqPxTBLjQQGJlsI7+/udCIRJGHAzVSOGOJGbVQGWCES13xNECDHWwh2RQEwiwc1VbRxHDixBOu4AEFEMwVRL0YsXLwIOEYVkyOJieufNl3/8/Vd/ff2rGzvLMlkWYu5TnXD33b3dmLp+sXFwcLCzsxNCMHc96WK69m4+fD2rmvv6aY+IGCCfoniOZA0ehoHNxdjzQ9v8RndDtSRxI1AI0d3LOB5ZCM6p2nU6gulRFZaeA7/sZ4RnLXKzcfZpB2TjkVMPqsn0+cS/dOZ6Yfvi66+/8tb33ty+sP3ZZ59fu/bJl59/OWRzZytGEIB9slh3chQzuNnhQrT+RjQZcbga3IgZxESkRd0NxA4QwUuBmRUFgZiMGHOW8nTLIkyzo/RcIq1r9flo/TOBGBBwlPj/s/dmMZJl23ne/6+19zkRmTX2PHdXD3fiJUyQlChbpmDJICQTJiTLgB4EyK8EbMAvhmA/GAb9YEOGYRjwLNqAAdmCZF8YEkRLtCFTvCIIWTJBg/S9vH2nnqr79ljdNWRlZsQ5e63lh30icqrKyq6u6q7q2h+6s2I4ceY4cfa/1/7/LnWrvI3aDU8GzM09SJEaJA10wj6pJqogJ+mydFlTYlbkxL6TpKKCvs9dSkklJ80pqWrOWQiz0dwZYalfLLbBCLfFDlNefPvb377Lx7HRaDQa9y5NgG40Go0HkZ//1V//v/6rXx1s83wet3Z3ZWOWZ3M4NIIMhAMiFIh4BMJVlZRwuBuEKyOLKccP4R4opSyXi+Q596k2sRBBIZ0R0XddzpmqY7EhMOvnLzz96M98/cVr28tr13fNwuuYUe6JuXXm29s7KV07e+bc7u5iZ3c3qTrCPNYuGfs2a/1sPQYV60pmkgLKSt6OiKkiafrYNGRVSEeEB8k61HXS36fJKKJd1xEwM5jtW4Gm01UOxcEdv0/uRZ+ExrG087zRaHwpWY9tWodMCBBgpKSPPvLwN7/5U48//phHvPHWxffe+2Dr2nWkHnCzABQQkDUPkEC4hTtFV2bQU7Lo+q4jzOAOARWUGlkoFMUqTDQCdXZ7hhokfXIqE1EAMEYU9wg3HLgb2YOAgImSNWlKhMM93N0DQHUcU0IUSSUlTcRMZCbMqlmZk+QkOTEpc0JOVEFKknPqu5yTiiCllFJS0QiM41jGwc0BjLDtxXJweOG8l93lrQNQG41Go/ElpgnQjUaj8YAyeHcmjQDGwZY6dBsbuTMpRYGUtNb+5pxqY4lkeFh4IOBwNxVRYQDmNprVUuON+Wwd9aciQpTlgIi+64ZhXCzHruvHcRisiOPR0/Of+8bLP3rt7XffvzQ6Cumx9j8kVl6HEcNisXvt+tapU5unTp+6cuWKmVElpRSBUsb6gZSyu7u7qtRqaIhQKCLVzSPcVVSlvotqwbGq7J705dXY1lqAtI4zDBGSrA02d3c3kGMZS21D7qmoX2It9YSaI2/04Gaf/RLvri8Th/oSmvrc+LS0c6Zxv7Cug5aaLRFhqnzkkYcvXHj+m9/8xjAOb11853vf/+HHn1wFEyDVuYKiEAHAiCnRYnpFAoBPuYOiK5E6IlRXUYFCkawqMoUW7o3CinA4hSmlKkUTK6uymsPBYha1i71mW0y/uSsxmhGkJJVZykIxs3AjXBBpMidDnySLpiRJNIlmiY7siSzIiZqYBEnYJRGFAHCXQBZh0MZYlqLJVW0SzomkSVMGeeXa9W2LiLi8VWad/OaPf/z5H9FGo9Fo3Ds0AbrRaDQeUH753/4v/9l/96vKGK0MA4Y8zFNGmLgJwhERrkwUAeCThltrcRilhKqqUkUco1v1hg5HHVvqNsX2uZXwUMFqyKcBoUCMy9N9f+HJh19+5tH3Pvrk+ntbNsnPKxOM1WP3WA7LK1evpJw3NjZms5lHaEok3D0lrYXYVYCOiJQUgLvX1qBHFZrpU0U194vMU7jQyvdj/Qant0V0Cqwn4QDhAgEiqXZdV00/IprAUrmZoNxqZhuNxi1pV4nGvQJZO96cjK7vnnv+meeef/b06dM/+OEP33jjzUsffrxYjkwdJRGCoCQVCgCJYDj2qqm5f6Z7HtDr3nYgAPdIOYtw6vSOfWbRYSAcB/yjEbBaxxwRHjh0FxJ7oRcElJJElcKpV70oUV2tlUxAJ9KJZJUkkoVZmMksyGQSEbJWcSMYFoYaiWGqbsUQMCtaQhmPcxcAACAASURBVMQ9HOGBkJS7jTSUcn30AVwO1p+bLa4s7uIBazQajcb9QBOgG41G48FFGYPFknO1ncW2b5w6TSDC3Ccp1sMlBIFxHM2cAEUJtTIiXIiURIQhIiIePhSrWi3MDWEMt7FaE4qIqIKek+YkSy/z1HfzjW9cePLdj6688cH26L6utTzYbItxHC9fvtJ1fUop56wppZyHcbBSpNYc1VIlIUlVjYhSClXMvQxl8ltEmLublVKq/4aI7DUGV74csRokO721eh2OGlI4NQ5Fu643c3dzs0AcFE8eQIPj4zf2NnbFA7X3Pk9O3h/AI09veGLfhm74JbZNbzQa9ysrowu4A/AIz1lPn9p85ZUXn37mqeWwvPj222+++eZydzeYtetEM6mcFF4yIAhBAOFgrO4iJtsND3OvGYMUVs8voRSzYRxFhavoiVWpc/20mFuxsk5RBgCHlxJmERZeEGWffwiAWoiMajuWRJIowYjpvqxqylk1CxOQwUxmMBG12LkOcZu81MAgPTgUBwLhHiV5LS0otYbaFKRHmIcBMY4mhdvDWFRHH98//cyp5dZv/vi7n9NRbDQajca9ShOgG41G48Hl53/113/7v/4357ZbiLDx+vUtltF2rohMjTBRcQ+zAlA15dyJJIaa1XGjVFVMg0YdoKqiGmJ0ycysjF3SAIZxCIpo7vqZm3nx+azTLFD72vOPv//xte+98ZP3ri63Fg44yHXbKyb9192G7e0tVen7HuPSd6LrOrOys7OzuXkqpTyOpQrKpUy+zBEQkb7vPRwBUakx8dW1o7parwqiV0XR09DXuvXcZyldcV/9qfbRnXsghsUiwsH9GvSXVTw9ql3Gvte/rFvdWHPDQ/zZK9xbjXyj0fj8OWyaXLu03X09QOqppx//+te/8tzzz7iXV7/36sW33rl2bbufbzJ1knrRDAoibCxeR3FFTdGIAPzw9TKijsmqFcuBIFTEI6zY7jBE+KqceW+lIry6kQGyujHCFEXoTvi0FXFgY9amYArJmlSVHuHBiCyaRTuRTjQJBawiOskAPTCGeNAhqCsTHjEGAggVqBDwNCKPQxSje1IRghJBB5wqs9PnBhsHcIxxHOKsvXW1f/4OH7pGo9Fo3Ic0AbrRaDQeaP70v/Xf/N5//m/MS1zXYWtYZiKWi1p9U9tfZlasdF0fKXkZgMRQD1Y7aBCiqkk9gqRqAkChR3YvpYxwjfBhHCX3QQxD1KKgsNHdgovHz22+9OyjLz39yKJ8vLvYdjCi2ihi7Y8RiHBb7G6TAE7XSpvJH3EyQqSZmdkq3gdT7CBBEffJfzGmemWfPJ0n4bk2+hwr+421p8b07vRwrUP7+lVVTSkXHfdJ2A8CRwMG75L6/AAWkt+n3IaC/OB8XxqNxr3JYQF6nRBIIiXd2Nx47vlnv/aNr25szj94/8M/+t733n/vg92dRZ5tCpWQCMLd3ctY3IwAIySC1cfs8MLqbcSkHlel2UT24iYi4PUdkJxCMcJRVWt6gIipShoBwhHO6Y4lcHAoVq2AVlKFSgIuhEL6lLNIEiaK1prvYM33oKHU2z8BhXV94RHhgAOhyqQUIIllNfFIpEAgIQjNBFVyoso4WiGWC+++9rpfOv/t337jbh7HRqPRaNwfNAG60Wg0HnS6ErvJS/FxKDNGn2bwxeQCHRFuQHRdIrm9ve0miJQk1YAcd9eU+llP0iKWw0CQ5M5ihwiE78QYYREx3zxD88uXdzc3Njbn852t7WEY3H3j4aeefvTcT33lhY+vDh9/sj1EGFYNtTp0VRSIMBuWS3dPqrnvRXU5LFXTxuZmKWUcR1LHcTSzrusAmE8R71zVDLmZ25QhqJr6vqu10iRruGB4kFNo4dqBpFY8V8F6CioEZGqjeq0B15TDw8qDYAUdRx40vsQcVmeO5VNp0Efr6Pd3abSC6Eaj8YWwd/GZzbpnnn3y5ZdffOH55z689NHrb7753e99b7lbzMU50hB0D7hZFIOvVeBghABHBeg11WWjit3GqRxacxJVN8PKBwxEDTBEcM99Y4oijL0lIuBYjdjaC9AgIERWKiCIiFBhJ2nW9wlkLdOOAFDcwh1eXaXdvXhEMKqxmVKEEAboqjQlEVkEKc9zP+u7ed+JQhPns0QV5rw0i7HUJMfFexdmTzb1udFoNBpAE6AbjUaj8c/91f/pn/wXf2Vz4/y1jz8aIEmSUGkLwADXLCrioFtYwCMYZkEGEdXIgsNQxjKOxUazWgrd5Vz12pyFFCC2t3ZAAbm8vl12dksZHRGU7etbanzpyYdff2j+3ru4vMTCY1ypzwK679Uju9nuYuGB3HUiDHM3s1I8gtRSipmJSATGcfBVkfK6KkjI6tMowljVULsHySQKrU9dRGoufa11JlgHwNYG4Z4tIoAIV6sNvmrPsa/J+UApaNynUd5QPbwNz99j9uR9XRN9e/7Ld5Z7TeHlzR/gHlvVxu1xBw9iOx8at8FJLykElOzn+ZHHzv/0T3/jyScf310uX3v9rYvvvFssutlmQAeLKFZvDMID7qtZThq0YcoxnIqXp1sHCjndkKwjBmM1aKsWQbtjVYU9xR+rThmDJNcpGe5uA9xiErp95Vi2kp4BJbNIVhWAESoUCsixWIEjLMwRHuEKSnWvjlrUjSQUCgkVSSpJJStzYs3wqEYcWZhT7nLuclJFSsxdDmBE7I4FoIx2+aHnZrtXf+Nbd/JANhqNRuP+pQnQjUaj0UDXz7e3r40ZMcbCo9dOI+BL1SQqomrhHi45g0QQoFnAoVkCHMeyHMaxlOI+mgGIIDzcymzWqwoQw7gLxGw2K25uRpEQCcpOuWrsnj5/6rlHT7/z0Mbuh4vBvUbxTHpvrNt2dI9huRQRVSWk+jRLbZRNOYQCoMrXtfRZSHcA1SFERTTCAdSJqxGHyBRI6O5mFgCEIhruAETE3d19nXOIujwg3N0V9YPFrJSIlSHjPafx3T1uJpWuRefb1lKP2YFfbg36c9i6++j8vI9WtdFo3LMc7Qc9kl4QQVKU586dfvbZJ1955aXZfOOjSx+//vqbH37wce7mKc0tOOwuq/jMCDIo6/rkqZ4ZAEjhVAgdYL3LkGq4sb82eh02SAERVfitFmFTXiGjjriaer4dPsUqRxjW/hsr6XktQCdKElGSEQzUzOVAjFYiPMLCLcwiPJNZRCFCirB+MKsImZQ5aVbJmbOsXdKcNKcaVEjNqUZD18BFVXVJw3IxuA+B3UVe/uQinn7ubh3PRqPRaNxvNAG60Wg0Gvj5X/31//M//dfUCJHBvadInsdg3XyuSRAhERKROoTTC8ZxNB+KDTYUkG5O1S6lDKZxdPOc8jgMw3IspawiDQOIYRhUVVUZKMO4HMsQ1H5z82z/0rOPXr6+eP/qWwsbSQ7uAEXozlU0YASi+mOoSkqp7/tTp04BcI/iUeVjMwO4sSG1zHltrVhKqRq1ahcRpYw557XhI8CUEgAPXw6Du1fNGjVTURU6mSXWOqPaFIRQXESkpgQtd3dtGtJ623rZbVQKf+EcMmo4uvK3tznHf+qG7352ybtxe3zGM/boIWv2341G4w5yQ4+s/WN3IAJ3C0Iknn7mqa997avnH374gw8/+sEPfvyTt99d7A7nH3p06/ruuBwpqgKu+rElUO80gOlWZzV3CuDuxTyntO7zXvWYs0Y5Tyo4J92Zq/sLcyvu9Q7KzMO93tF4FLMS6/jB1eZhtTECCJhICYRZgF6Hbu27oFZ/MxEiQskkkkV71U4kT9XN2uukOCdGUuQEJZKgz9p1mnPqZ33Xz7q+H8ZhGEeIFOhye9uFZvH3fvCDrz788A9+9O07ehwbjUajcR/TBOhGo9FoAMCf/at/5zt/909c+uGzQNKs8/lmLHW+OZtk3Kj+G1TpRVIEl8vlsFwSYWZlGCgUgmBtIyXV5XKZUlIVDx/GEREUiAoID5h78bCAmcWwO2xfPdPLEw9tnt/UnWEoBdVC0WpUD7DO2HH3YbncEZnPN0heuXJlY2Mj504Eq5rmKTGwJiKWUlR1HW3vHrUEKSWthc+qWkVtEZ2CDQF3p1Aoe3OsM51ygzCNpa1xhKu8QyvF3cPsMxyH+0t6Pp7PXwh+MP1P7gU+e5Hy8WdLK4K+LyHw5OZGoiRhEsmrB53IRk6nUj6V02bOmymdynme9L/9o1ffvr79Ra9148vEoevGMReZqfd4Pu8ffuTshQsvPPXU07u7i4sX3/n+93907foOoGW0CFAkSR15JaIi1SvMzFcCNFf1yDVtkBGSQlWFIsL6Yr2xmbrA960B1uETViXtMI/wcLdq9+G1bNnthhbT65dUoCIKshZS1zVDXetaY01lCCFAFukomZy+oYwkyIhO2SXpsiR6EnSddio5SZ81JVFl36WchHAlRGVwvbq7s+1hRvf45y888X+/8f5tHrdGo9FofBlpAnSj0Wg0Jk49cu2bf/5bv/uf/WUq86xLfcpZqwBtAQ2Ys+83u24jdbNiZRgGK+M4LIbFLhECKKb2TCCWy2G+uaGqpZSd3R03hzB3ubiP42jDIKI5BUsJj3H32kbuHju38dSjG1vLsn1lIBgIjyrmxpTAE0D4MCyLWUrJ3JbLJYCNzam2h6SqrOqgEynVeSPnrKpmXspY653JHBEiTCnVt6YiJEFOqTpZT8XaNaVwSjWcWo51lG7NrAeQA+6ed3MZR7fVOu+1dR8Q7eyGdaz3vpnv57lWJ1Tkj1dj70hF+R3vG7gjGvT+uaEVs9/v/AtPPP6XX3nphBP/r6+93tTnxl3gpJe+CKQsZ8+ffuWrL75w4fkzp8+++fY7r7325htvXtTc5ZS3t3eDkiRVg7B1pzcDhMg+AZorCbqUAjIlxcr4C6ty6TpCy2Pq2GY1EIuodc6llFql7OFRQwKBGhKIMIQfvdyui6BJSvXfgMCCqKsrnIq2IaQKlVRCyV6ko6SgIhRQhEZouIQomMgkkRP7pH2X+pxyViGqAYiVsYxD8TDJu+N4dbEszjG8y/HMuVN35gA2Go1G48tCE6AbjUajMfHCn/zeH/ytf3GZgqNxe/v0xkZZDkIkFfMoFsvRhsG6buz7kSokulmXsqasSYRAjLVd5AC0m/VWrBQQZ88/ZGHu7uFUATgMQ7gTsFLKWMo4Fu3nZx4Z02n83o8+ufLaiIijDcV9GpeZz2azs2fOiIiZqdZanyl4UFXrkNau6yJiGEZgdDczj/D6Vkx4rUIaRxOhqg5lnGqiVUiGx3psLFY1SrW0ae3kGOZWStWsrZRArAKBcBNLis9fVrvb5h4388T4tEu8N0XqO8UNh4HfbMo7y6FjcXuBkMeft3ewx6UVs9/3ZJFffu7ZE078T97/4B+/24olG3ebPZH24CUxAFB47vzmiy899wt/4hfOnD5/6fKVP/jD77z99nuBpNIBshxNE0EvxdeeG9x3X8BpVuv+8nB31ldEKSLg+h6ifmrvPqKalXlMr6/LqLkymHYLM/jK93lKJoz910gCJITUSV4WSggorI7UKy+zqGkXdRHhmlylRmeoiCKysk+aJRI9SfQ59VlzUgbGsZRSSJCxtbMzmluEUSPPr5eyDBaO3alig3zr/3nt7hzERqPRaNyvNAG60Wg0GhMkfuuvndPFe376id1h6LsuShEfktId5mElMI6+XAw7W7nvu9lM5zNNEuhUFB4W5m6IyKqK0DArI4CUk7t5WETUyMAuJwJCKaXYWEopxtRtqM5Of/zJ9nvvX3rzyvbW0o0S4TdQcN2H5SIl7ft+sViYmeYM7MnDNXenFhyZ2Z4/I+DmIEQU1ZyxjCIC0MxFqCpjMQ+PAIUE3E0oFK1LXs083AxTqg9YvTgAUdWkbvQpm/5Bk89uWfJ8vIL5oO2u+45Wktw4KX/m6afO9d1Jpnz92tb/8uPX7/b6NB5U9ne+cvV3/WD6TSehCU8+9fiFF194+plnPvn42ttv/+StN9++evV60l6YA+IRdA+gjObu1YALgb3EiFhZb6zU5fqXCEiQ4que7/XK1QkAQAQEvN4jTet8YDp3uKGWQmNP8F4L6QSETMJEraZorHcxUxgG1oqzwDVCCQGESMqM6MhOJCfPwj7LLGsWJKViCuIwD6uienVHI3YWi8GMOetsNuyOu3AjF9p1I3JX7vyRbDQajcZ9ThOgG41Go7GHLK6P585iOYRj+/p2IjHsJDEPAlQRjFHMF8NytnmK584ndUkdmYrDnSXoIQS6bsbwsJJTdrdipdY755TMio2jrvyXERBq188Hcw05c3bj41eeuPTxR9vfeXsYFoNo2acdT0RE2O7OdiljKWV3d9fMUkoR4R6OGhE4tTBXVc4OQFNS1TKOIDXlauJcSomV4Uadu1ePjjoetqbPc+8pUaeMUoqKUKRumpAERSTnbsQYFodXe4/PR8K7YcnzSUqSP2Ot9DEfbE6+XwKaBt24NZs5/dIzT51kyivD8N+/+v1y06tlo/FZONohKvsE6Jo2HKoqwtzx+Reef+HChdls46NLb7z22huXPrw0FuTZqQARENKmuOMCn8y46lI4FSvvX6jXcmfWJInJIkxrjzg8Vh/CykAMAANBFUkS7nv3MB7hAXesB2ABoB/YygBJFcmiCaIU+JR1aFbMioXVkVmCSAwhRZlFsmCmmCf2ypyYk3TKPuksa1IhYG5Wxoigptr7PoxjcbfA7mIslKx9z27XFiXJODqsDF33N7/947txOBuNRqNxX9ME6Eaj0Wjs8ad/7dv/+1//1688JY/8eLhS/FSSTtRtjCApiBC6aGzOOvdy/erlxXLhkkeX+eaplGceVBWBLJajCoRShiHgqlqHmnqJ8CBk8la2AEKEmhIVyQHYS08/sfuzeP3dK5e3dooVOVRIPI0inXwXx3Hc2NjIOddowQhwSvqR/WVGVYWuqYPVXoMitcG2tnhWnSIHzR2kJq1hQWYFoKyHwdYZupuZTA7RRkDAcISbWRGRcWApJcLjXqmDbrrh58b+Urt7ijvVAXAvnM+Ne5o/++wz83TrVsbo/uvf+/61YfwcVqnxYFMvyGv1uRpeEHDAI+LRxx596SsvvPKVr8zmG6+9/sZ3/+h7P/rxa0tzD4nlsDYEm37TPVBtMlaSMyhr+XmaEvX2RvbfZoQ7yaTKXPus99kbCQGERx1RRZFaHC1gwM3LZP18DBHwIIIEI4DiAUeEGxGdMKWcU+pUs7AT9sJe2Al6kU6ZFUmZVJIwqUA0KAEEhaQHx2UZxnEcB0dYuDugIl2STkezAWHG3XH8YGvnn731wR07bo1Go9H4EtEE6Eaj0WgcYOe8PKsfXI1Hogy7hdJ3w86iSsZZdYwCuKa0HMtiMOm2C3Qwzk9t524WVJWUqAoKQhDuhvDquZFUGAHWEaZWjSvcHCTE3QEPwh8+s/HVF57+2oWnPrm+2H7/avVsPqx4ESDDYxyGjfl8NpuRUv09+tmMqhFxqKW21qPJOpjVOVl0SDXoUK1lSrRwVgEaCI9iBevWZ21Jmnu4u4sICXefIhLN3cws1QYnQLPRpkzCz59bRgIehSv/yntQPL1f2G8qeg/uxlaE3rjrPNT3f+rJJ04y5d/+8etvbV2/2+vTaKx1572UPnLlfRFdnx997JFvfOPrjz72+DCOP/zha2+99fbHn1yB5hApbtMAJ65MLfRAjzRBqpJHfnA5BUiQ4m7hEeaiIioyjbg6IECzauHuHut/nQx3rNTnm169CRAUQIIC1FBockoeVDJL6rtu1uUupSyShR2ZiSzIwkSIhAhVSIFTSogHI2DmdET4MIzLcRjGAXUvCDdns/mZU0bZKWOIlrC/9903vvrYuTt53BqNRqPxJaIJ0I1Go9E4wF/6S9/60e98/U/8xd/5B//hXxhpW9tbu59cyUm7nPt+trvYGW3IXTeOZbkcmbIFhxL2wfsGOhXOrOmh02d9HJe7u/PNubtd3956/NHHzp45q6opiQiLF1HNKZdiQMgwuhkDOSVqnJqlX/jZn94a9fX3fk8IqcE8e427gEcQBnfDWEoupb6tSfv5nOSwXELXw2yxihksZtb3NZZwqHXTpVitfRaRqisLhcKpMSnQ0OrjKKhT0SXWuT+1LRvu4W4sNsXMU1RFdLGAH7UQuSl3XLK8Yf7hSaY/uUa5f51vlkN46MGXkhtu+70m9Z7w6H8h3KnT44R5iY27yL/6wnN55Vl0DL/1k3f/6Qcffg7r03jg4b7a58kxi6QKPUISzp0/9eTTjz377NNJ87vvfvjqqz+6cvV66nrRZI7iTkmqqikp60gp3fthCwiYcpKD57wQFJgZJk8vQXgZC2vlM6eBWb43PVmtnut/bqUUKxZugbLy37hBNjNWW5UoGaJgAhIjCfuU5jlLRAJykqo+C5jIRKQpphBZVUWCEYgxas3AVEjtZuMw1tiLcRwCABURWWRj3j328Jlzjz9ybXt7cXXXS9gw/Lknzv8f71++ewey0Wg0Gvc1TYBuNBqNxmFe/sVX/+Bv/0K3m8d+d7TIm2eV8PDBzMDiMiwGBCGdO90jPEhhhI2DmRt1GwyzcTkEPCLG5Xj16rVhOYLMOaWsHq6qKWVzEyLnhPAwg3tIN0r/yKn+uUdPP/PQ7NL2eG1pfliDZh3uGhHLxVJVT58+A4Ckm9XCZoDuYaunOec6QW0l5pzrBLUKai/RfpX/4+axjhxEwGFhZravlnqdd7jOlXe4B4KkiGpKqsmk1LCiE5sv318crz7v53h5+p61rbgl95rKfJSTrOEXvhV3qvfl6Al5P55U9zFPb2788cceveVkr16+8nffeOtzWJ9G4+BFgADcg/QgEGWW+5dffvHCC89vzjdee/3iD3/42uVPriJkY2MTFA9YxNr4C6jRgO5T7h8BOGK5XNZZr7ubyagDpLDqAq/OXeGOCJIH5GROc1/lGlZxOlBvsNxvJj1PBAAk0U5SpmRhp8zkLKVZ36mHhCeCHjaWGnrogFOEEMRY73mmiMPwqG4eVFFEmI0qSMpUCxG6PJv1s3k3n+czZzdSSkMxJsrIn/mDN99/opU/NxqNRuOmNAG60Wg0Goch8Q//3edKXkS4Qfo+z/pZDEuiMGXtbLlcinYp9W5ezLKbpOwRy3FpxcKDCICatJb3dKkfluNyOXpEyinnREJUkyoYqtJ3qYq+ZViCCXnj9Pz8Mw9tfu2Zh//o4ic7y90CSJV5qwf0arBrkMMwaEpnzwoAM9vd2V1l/tDdx3GsyT91PKu5x+CYIuXH8ABQh7sSqLVNoATgVpt8FGFVqN3dzd1tnVC/yg2aWqERwbqCQQA1ZVFUPWrt0gPofnBL7e8L3y2fUff8Yg/ol+x0ujdNSxqfjj//wvO3PIof7S7+x+//0FvwYONzIvaVP9ffHI+IgM/n/aOPPfqVV1558vHHx2F8/bU3f/TD17ev72rKKWUPkhBEVCnYvMrCAGs/dDV+DkQpFu6MQ53NK5WaEivrrrCVlTMFInvjtGS6i5iekpxue7xq1li7fhzqrg0QUDKJ5pQTmFWSMpGSlKKAw8PCixV4MIIRCiirWUf1sw6HO6tpWjCokGqcRjgpOaXNjX7e9/NZf/rMqdnGrJ/n3OUr29cXgdBU/Po7Lz75zOvv3d0j2Wg0Go37mSZANxqNRuMG/NJ/8q2//x/8KxSoJuZ+8/SZWc4JRVRAltEpWTSbhVX5NgJ00s2sDGVcDuNiHIexlgmJyM5idzkOAgR8OY4EkjqSd10W0qyoMCXpu02RRM3O8vwjp37x577x8fXvvH9lV1bmxAEGpwYTQEYEoozD9evXzXwYxgivdc418SfcKUoCVkAJUZjVCcIMESBRm6JSq5/3tQnDp5j7ydO5Ng5dNJES4VV5njwe9x5DWO2tDYSoiIlzSixa7eCbOTbcWQHumLmdvHL55Mv6VLM6XJL2abizutWhuVVr0C9cGjvpCtxsvxOM42ZyB8+0e7NnpWnZXwCvnD3zUw+dP36ahdlf/973t0v5fFapcc+w51uFk14yjtoqHzv1kaexCgNcWXAADDBEAuHu5cWXvvJzP/czL774opu99uM33nrz7Q8/+Hi0EHFwqFmD6/lGrBKNI1bpyLJ6y+GOALB6iwSIcIpAUtWdYzUXAIDDAlRQAIStM5Zr57eg9pRbCbcpNDFiXQm9/o0SQMlONJMa0+1HcYKw0Yax0APhCI9a4uwh4YxQhAL1rxBCipJKUc5meXNj3qn2SWdd6tL0oOZ7SOyGhTsvbw8fbV3fLdz1Qbr51fP4H050WBuNRqPxgNIE6Eaj0WjcGAoCqoAJndFtbvYoKiQEMwYV0ICsWmQOhirczUopo5XRbTSz4h4InBqHYRyLu3mN6ivhDnhxGxeD2dB1OamEmWpSTcUkTJ44f+rCUw9fur578dJWcXeyYE+nZUQdsmqlbG9viyghoESEFdOUBDJGQZWEoRQBNQhUy5BaECWCdfkzScoUQh9RvR6n1iYhoiQifMq7j1qNzelvHaG7/t/DuJKkwVLGUspBW4C7rdkdFeBuKMkdXZM7pU1/2gjEe4T7ZT0njj1IN1enTzrlLeFn+/jRWX0q7kHh+4HmL1x4/vgJAvgbP/jRezs7n8/6NO4lpqvE3fvSHrx2M/ZeIyigIryaT4Do+nzmzPkXLjz3woXnu9y9/d7b3/nOH33w4aXdxRJQ0lGNv6aZrSMlaonzSkTmepmx2sSYNOhV/GAdUwUhYl/y4R5rZbx6ftURVLUPNBA1htlXS+D6n2n6mGahERJRPdGMMEZhSEAxWYQJiXCGS4CEqGSRrJJFqgadVDRLSqKJs77bmM+SsE8677ouaafSZwHMwxyg6mDxybWtbYuFY2t7o8vj//b7r9/R49loNBqNLxtNgG40Go3GjfnlX/vNv/9rvzIievfFWDxcksKdiCTqERaWUpViUctuVOnByMoNrSM73cxGG4tRxCMWy9HcrGQ/xAAAIABJREFUzGwYFsOwXI6L3d2dYTkuFwt3F+Huzo6IpJSHwZA3+o1zLz/36NYwfnJtZ2eIEijVqXlVKVS9Psxsd3d7Ptuczfuk6u7FbGNzkyqL5ZKkCDUlrtVkn1qJ1Z2jbm+q8YhkOMzczLq+V1UrxcwiIudM0t0t7IALNPYG0a4cORDuY1FNqmUUkVigxi3uayMfo/x+dvZMQg6+csN6spst91Otz2SmQR5a4uEZRq06B460w49OfrLJ7izk5AX+xRdB3yb7qvW57yhMJ8OhnTrJHVi/c/uL/UyfvpMzuSvc+Gy46TlST6KVM8/eETl4AL6QM/yu8bOPPPzC6dPHT/MP3nr7Dz/+5PNZn8a9x6f+gn/a78Y+Z2auL+OEQBWiMEQYopC6cWr+/IXnnn3+2fMPnb986ZM33rz4nT96dbH0ACOCXl0yphWOkPWXenUZ5coX+uBGVZOOcIpQVYRTajJ1tYYHhqbQq5CM6lwWXJVQr7v2a81zrK/Ue9durkRvRjCMMBLh4eEBC7iAmcopl0IEEDAruyRdShtdP8+pT0nhwsiqqZOUJSfJKWVVFWTVLuVOJavkBA8UgwPGdPna9W3DwmO2nc+oXxvzpzxWjUaj0XjgaAJ0o9FoNG6KA4+9ePny248VG65sXZXZPFlROFIKhAfomcKICIJCSopAeJRVgJ9QUtau70EJyOamFCvmFvAqjo3jOCwWi90dUZIsY3HAAsuhDMZl6MsXNkek996/9PalrU92xklGXVX+cP3EsVwu3Hy2sbExn5/d2JCkonrm7Nl1wRImFwxGeJhPTTKRqi+vS5kBqU24nLOIeEpTRCGBgKpqqMfKCnIVGYSAmdVMe67aixbuHiBVNedcyjilCR3HpxpzfPwcjtGCj3n9duSwvUb4+kEcfLr/CQ+q4fuL1tYrsToih3XRlaZwvHZ+ZGX2NupgxdqRT6wnY+3d2F/2do+xlkKmIv3V3l29uzdl4NDePnxU9rbu4MH4Yrb6llXbJ61SjyMfuxk3nh333jlueTd4b98nsT6ReXgFjtX8V6P17w+E/JUXnjt+mj+49PFvXnz781mfxoMLQRFKdYsgKJoSqaCEl3CBs+/z+YfOvvDCcw+dP7dcLP/wO9/9/muvL0vk+UYKWS4HEaFIvbUBYcWqn1hKqklVFJMLWB30tLfwyZIsVprv5Oy8enevgHq1snvJEZNYbqWYFSsl3GEG+KHrwP6LNYEMdGBHSeESoUEhhYlAEmZVMoRUUQGU0Sk71V61z9In9glKqlAVmqCZKvU/FZLBsBjMR1hECYQJRs2L5fUt85EktPS2udS/+fu/f/cOaaPRaDS+HDQButFoNBo35Vd+7Td+9Dtf/+N/5Xf/0X/8F7dK5NEy6TtXs0CUEKpqkFOmu2ruu2kMaIAUFU2aVZNoEsmiiYQqRYSqFKHIrO/Gvuv7XEerRsAiLDB6DBbLEuce6nLutq5d53df337rwwBs5el4CDOLGHTMPpupSCklIlLONX7Q3QmQIkJ3esRU71yrjNzXKxBhta6pjJNLaY2kd/PVU0SEw/e0ZyAiSinVMzrCEREI9wiApKhqSu5uEceKSp/dG+GLrSE9Zukr1XmtPnOfhrx/EPMh3W5F3OjF4xd5YHYn/ggPCZf7NOj10m9e+XonfEv2acUHymYP1jPvvc5Dyv6BKdcbc6Bo/9AumGT9e6EA+WY78FDHwa3383q6Y/obbpvDO/zonpuWF/tPwL01+Yzl5vcef/KJxx+bz4+Z4N3tnb/xwx/fN4J6415k/QW6SdfpqhdZRKkK0RChasodhQTGwUU1af/k4489//yzTzzxWCnlrbfffu3Nty59clVyn7oekKBU76yoY3oCql4vxSIiKkm19vpVfbneSNSVqNETU+clq0NHjTL2lW/HkR+Jen0m1tcGYnJtvtkPSgAMEEhAR5mJzCQlMBMZmkSUstKRKQwCQhGEILKgU+lUe5VepVNmVVWKOKvkjAj34oVgjV+smniEsUs63xiTb5dSRAdx6eYZy19v6nOj0Wg0TkAToBuNRqNxHC//4qvf+Tu/4Kpl3P14uWApy8sfpChdl3KXADjCIoIiOad+VptFItJ1/aybJ80BmsdstpFz55hqgmIl44LhbqUUFRWRCJLMSfqcIQlIKXePnDt7/uy5re3x4jsf0jEAY4QdNLOgqAcCLGbL5XJbdWexS5HNcfRqPG2mqiklUQ3zMo6qWi013B21YSkiIuNoBFNKi8WiWMk5V5HazLgagLtWkadKbxCAmYlQVUspZgZAqqhdjT4CZubhYfublCcRZE6uQd9S1brteupbfHBPEjgiDhzWTKcX48DL+95bKa5Tk35/236v2nef6HpUYTygUty4XPrAJ264hvvX7ZD2faCa+tg9c1OlZG1DcnjF9u2NtRnIaiv2XlxvQBzMtdz39PgVuAHrHT49XR2IE378znD8aXbSszdu9vToDHjwBOTBQxIADu/SaU48eNIdnfNxS70xsffPfabTJvJPPfnE9njTXMEaPLg0+zzXqnF/c7Sz8bgxPZPiWzuPRZSaonZ3q6acSIYbwlR56tTmV776yisvv3T29OZbF9/5/g9e++DDj4thY/NMeADcmOdSirunpO4REV3XiQiA2rF9eNl7wYSxSmWeuqXdQ0SSajGrNxu1x3vaPgLOaX5TvjJQ1Wc3hN8gSnZ1jWJAgET2IrPUbeS+E+lEkmgWTaJJhQyGV+tnBOoDhqNe16pHNSXnnJMEzGERYe5mXspQAzaG5XK5uzOOS0mST232xWO+UZI6y/jkT8nWpf/5H/3Tz3KcG41Go/Hg0AToRqPRaBwHiX/4156T69eQuGOSinWnz8u4rQLVNAyDiG70M6uKjNNRTTiwu727e2035UzSAlf8cpCimlQpGEupA1QBDwQiVJPUIZ8ACZHaMlKR7MxnNH3t+Yc++Pi5/+/HH1zZXYbAA5PPBzgFxAPwKOM4iKiIigZxbWurVh6RqCXPAN3MxpJzAlhKqaoxKauRs1MoUG2CDsNACkipFo37ClKrLwdFgGrugQA8gjWvcCplAkkDKD45fvg6UGjNfjX2prWUn4E7WAZ6kznEvrrOAwL7Dbbz1oL6Pp+Nld12rD842U2s5nxQyT6wrENa4r4pj1urfcrhTavPDj66hQZ949fj1tNgn9Bc5ZjYp6ff8IM31V5v9PSGyvtqm+JI18DRk+gkJ9WhhXwqS4w48fRHF3Syt262g/YfnRtWK9+y1P3TC9D3LyXiP/p//+CLXovGl4C1ncWe1/INpjn0+EB3HAP0CJjDIYIwDLaAm9sY8NPnzr3y8oWXLlx45KGHPvzww7cvvnPx4sXFcjTHYjG4OyIYNPdwH4R1nJOoTN3M7tNyYp9J9EpuXv9crf+vrl8mMhl5idRJER4kKMDUybX6zQuEh3sdR7Wa076OxlW/YBLpyAxmTVmTipDiIR5agh5wDyFFUoR5ICYB3MJMhDl5rzZT7VVle0lYeDGvMjlUJeckgpx0Nu+6XpJsntrozj351Ch458pOsbiymM8uveuPPHUnjnuj0Wg0HgiaAN1oNBqNW/BL/963/vG/84tnt3beffRRI1KXuv60hCVKhJBUyeHuIKkRXh0vymDjMKacRSSI5WJwj9RnICKsmJFMmiIMhFBEVESIEATDuSrQUclIs+hOPXGue+W5Ry6+/8nOOJitmmUApqGukzzsxUYZVXXz9OkAdrevryqbGUA14pjaYWYE3UyYVv4b4e6qAoRXu2eVKkmLqoqg2jFO7dxVxahKLYGSVeq9cDWYtk7uXhvTyX0qlnK/kbxX+VSi2z3GPidiYFVberjpzBvK4YcqeQ/O44AR86EJcGQfHSNJ40iR66HJbvrWuudhfzn2XT066911RGrf//gG7s1721krePeVmx84syZ/mDg4/XEBjDfoH7nlHoiDPQ4n7wtZdwecfPqbHZFj3joBh87q/a8Dn2nOjUZjYp+UPJkbA4e15tUF6kY/HVFfr7+7HgxDzQ6UsMEiCnw8ff70U08+8fWvfe38+XPL5eLNNy9efOcnH39ymTqLEC/LiH3OWnsOW5juEDD9gGOy0gpQgAO2WqueZ65zYIOYdO11zgRBlyCnzq3Vtbfq0O4ebvDVIlBdog+MvxEyUzLZgan2gXtYuCNcpmREIZJI0mRe3C3MzYt5MQ8lU8RgMUh0GhIGLzDzMI+IwGzW5blqktmsO3NqIyvmnZw/s3H6sccuXbk6W447O8vNbrF9Db/x29+6QydAo9FoNL78NAG60Wg0Grdmc2vn8tlN5oX4nKr9fIPjKB6bm6eHYXnt2rWxuKS00Z1CqLvZOERESklEVEVVGYiIbtZv7+4sFsvcdSqElwgPMEgPRyllHOguNRA+DO4pZUfatktl1LNzefScXF1wa2sK+5tqkj2gXJccmXkp1nWd5jRamc1nXdfVwaTunlKOCBsLpppdqqaUVCdXx6jqNik5JQqrPbRQAFAEQjdbKaG1hcm1K/WUBgcA8PBwczMP92SpaFIZVUiO42hmK4H26P6+pZ51G5rXbWtkn/KDR7XLwzJwHH3tBlPdaiVOvlqfSp6+xcwP1C1/HrLj3nDvT1Fye/DpsbXW++Z/dPobLXGlk+yb4JgVu6F2fJL9dqKjceynTv7WSWZ81+bcaHxpOZl/Dw/8A0xlxQdriVf/8OiXcX+32LoeuQq6XnvwvIyI0vX6/LPPfvOnvvHNb37z4sW3vv/qq7/3e79/deu6BWjhxWK0WFscyWTogZUKHfsvd1ViXq0qsCcucxpohdoTX2MnqkRcbyRqTbSKWITVuIgAIhiGCARr4sRKffajO0wABROYQAVgZuYDyur2Yx23EErNmgI+ZSPCgYBQakU3WTs4c5c77VWoSlWKcnNz4+yZMylx1qVTG/Mk3iWe2ux2zD/e3l5alM7eef/q737/3RMd4kaj0Wg0ADQButFoNBon4ed//fd/49f+JbFO1EcVzrrZ6TNc7s67rrc+9dkMAZGc3dGZezfWoZwpZRBuxk4C0JT6blYlXyLCrWq5EWQIANXEBCHCza0YhkAGkyadUR86m75y4fkdf//S9Y/KnjOvgBK+bh6Gu43jsLOzM9uYb2xspJSEdPekSTutns4lFdQGoexvuwbgqqytQg8XFwBmVrwAoAiVpVjU4bSrNuJay15nFdbcwjqWttY0TbI1KapiNg3IvX2OatC3bO3fbHFHfYOPn6DxALJfSr4jivDNTqq7oee2E7hxL3On/JG+aG4ercm9Auf18KADb0+sftT3/sa+jwLrvt49YuX7tFc2vZ52Gpgkgo35xkMPn/3qV7/y9FNPLZfLd975yetvXLx69fpoQc2AihJI1Vm5WiNzEqBBAFL9tGqP3d46rKepim7EygG6xlmQ62yJmAY/RZ2ZqIo7rQQi3N08DOEBX2cPHtrS1RIBhSSQEXX0iiNKwMHqCr3eBSREoLUIm0GhSFJl13V9zrMudSKZUGCetcsqwpQkJYpKyilrZEWSCBsMHJG2XT64/Mn24MXsb/3OD7/5wsM3PxUajUaj0bgBTYBuNBqNxon4lV/79m/++3/Ol/QuRiunTmdoiErHbr65Ec5iGEoVZoMIL6Nbybl3j8VikSOCoEhKfXEHEOERbsXNwr227iQIURGBWRnKYMMSklRz1hwF55N/9aXTl3fxxntXbVmseACowe22lsYi3EsZt7auBeLcQ+fd3cZiVnLOSVVFIiK0mn6QpJnZXkCQA1JNMooZAQpLMbNCkMIQerE6aW3n+sqUUYTwyWgxpneDgIhWrV1IsLqNaEiY7dV43Rb7NejbVp9xsILsGAeDxgPLoU6aO8INT6q7pMEdPcPb+dy4R7gbX67PHa59MTh93fZ94SY1dHp3/8RH54N9WvKeDL1vH0XEvqLg2Fvg9PHqcLF2SqaTzF16+JGHXnzp+ZcuXDh96tS7P3n3rYvvvPfBRx5CETKLJKEySzAoIKcAYawdM0T2CdB+4JeXIKiaiOleopiZm2pKmqYwC2EE3K1EoUiNu/BqylEdknzlzeUl3A/WPh/YVQIomSla/UUAVK9oUjjVRAsppJJJJSclgoSKqEpOujHrN/p+3udOJSHg3ifJSlGmJDWMw8LLuOvQEqOPwaSCzd3t3UvXd3a9yPbuv/zKU7/1o1b+3Gg0Go1PRxOgG41Go3FSwhhd4mDXU1l89Emf84ZgJsiqbgEmzTM6EJGUOuuEVE3uMZ/3qOU3KY1my6EM4yDClNNKgEYE3WMcR4qIcPSiw4Kqfe5VEig+FmRunJ1/cn3x4eWtH1z88KNrO8vJCQOxyvGZht86h8XuQmXY2DCzUgoYZjaOBYB7uFvOXUpJhKUUW7lqAHQPgKpaSgl30WnwbE019HAKVVImKQRhVQavA1oj3H0YxohISasArarVclqEbjYSIiKjLpfhZtWy40jUPQ759R46FDea5uQcbf7fcIa3tEFoKt4XQBI523Uz1U4kq2QRc1+aL92WZlvDOPgNRm3fFjc8vp+9WvOY0+YzlkVz36PYyKkXzSKdShZVUlb/EfCIElHcF2bXx3F7LPa5eKo07hGEPJPzma7rVTpREKP7aL41jtfGcTD7PFbicMnwze3X7xG4Twree7H6UE25gdVigjLZaEzjfvbLyOTJNnIK8d2/vDqz9RQBTL5XNQdCQaGQ1UA5EOEh8DNnzrzyyst/7I/93Gzef/D+B9/93qvvv//hOPp847Q53EOgpEB0lUDsgWkU1DRrc6yMNeL/Z+9Ng+VKsvOws2TeW1VvwfqwdKOBBnpDo7cZcmZIjiSKtIKkOOSI0jiCpBQKOxRUKBzhLcIhR0gO29GKkO2Q5OWHLP+QLYapsCWRY4q2htTIlEmPZVIWZ9Sz9N6NbnQ30ECjATwAb6uqezPPOf6R99b26r1X7+EB0zO8X3fgVd2bNzPvUpWV3/nyO6AVCV7lhkVAIKx+Wkgy3VKNZUiXo6LQTaqEEFkGzCBqKqZiWCUxBhHQaDGCjRLck+wzAWSELabMMCUhNFBMds+AHsk5cuycY5eSIRsAGCEwEYEhAopYDMgEBgYpYYcJITtSZW/MxqISJSKaiUkslb0Uca1flkghCLX4MWj9zkw3sUGDBg0aNBiiIaAbNGjQoMGs+MJ/9dWvvPinb0Or0y0JQ3CxJHShn3OaiDnO2moGZt6zZ/LMRC7Ryj7PnfMhmKiCCSEQoWP0zqtaCMrIgCiR06xTwYfoypBnPkMkFc1inDPAVifKCVXtdTf6/Z6UlgRRSeMDI0aNqlYWxdrKivOeCLUyVQSzKgkhEQPYCPVcQRQQkYAMzdBENS3itdowt5JbVbIuZEpTXU2NJ3vHpLFOFSY9WNoIgMRsBimvoakZiE2hhDcRE/fqjDGoYXb673tZkff9gnnvT8/PPTI/f2qus9RuH8yzee+3uYUGsFKWN7q9m/3+lfWNN+7cvdXv34d+Vc9Gznyy0wmqQVVSbs1BJKcW4iUt3noIayHcp6DFT5x6+HCrdSDLDmbZnHdzzrWc221LK2V5q9+/1S+urK9/sLZ+ZX0j7BuVP4Y55xzR1F0KtlaG/WroQJbtWMbAVnff4udPHC9Egmopknj8oKpmydZWLdkfVHcgMf5JUEpJTopYk4voCBNT5okGLxjRETqkiyurl9fXd33mW+BEp/30oYNnFxZOzc0ttVu0tWXERowfd3vXu93319Yvra591O3uVx/G8L2xtmREzjzupFFtqm0oBlTrUJCclgENHJNHjxjBpqSzw+2b1uZM+G9AHf6td1VZgxEBVZRQ5zrtM6dPnTl9+vDhIx9++OF7lz744P0rK3fXJSqQqlUZAgERUKDKKCwAaACa3DCqNKSDs1BTGXqApZNGqtZfVZS4VVkEqxh5fSZmCBFYTS1ZbVRsvCmoglqivlPoeqAorz4yZgTmANpE897niN7QARgogjEhAzkgJmJEBmQENDU1JCAi5vTTSmOUQBwcAJgAmBoRkBlqZFGO4phUYwjBOyICQHVzrY31fo8ogmKrr9H93ZcubfPENGjQoEGDBlPRENANGjRo0GAX6IF3UJTQx9IV/ZJCoLKbYUQAQAb2ogpomWPHzrFjZlULIc7PL/gsj1GTVQU5x0ymmOctMJBYuCzPvKfMmZmCMTvATFWJvYGVZTlnnFjuhbmlI4cOXLn8wfLt271SykpyVRkmjvCsHMp4Z/n2wcMHO3NtizYgqdOUkQhVtd/vM7Nz1YCY5M+10pkAUaMYISBEFQBIPo8Dno2IaoFzhDRnhTTJBFNFJAOQKIhAADGKqhKRalQ1ZEYVSH4k1bGDafRm3DtRsY1lx1ZEyGba+nuDMvmeBgI8urjw7OFDzx4+dGpubrfHHsyyg1n2JBxIW5b7/TfurvzBxzcura7tdzfhWLv9H3/q+VlK/+o7l/7FR9fvpa1t8LNnTm9F6c6OA1l2IMseW4QfOrYEAEH14srqq7fvvHTz1nrYN1IYAH7p6aeeOnhgq73/w2tvvHb7zr409O8+e+Hhuc72ZdZC+Cv/6hu7rfkXHjt77xd8FvzKWxfvnYA+kGU/cvzYDx8/ttRuzXjInHPnFhfOLS58/sRxALhdFOlJeGdl9R47M4kqpvnJwYBi3rxlSDxX5hHV/tqqAqp9UHHKFTWbAsTj6xPGWxgJAo/Hg23T2iCbIhInqkqaJocM8h4ATMrM+8MHFy6cf/KhkyfLMl66dPmtty7duL4cRVQtSG/EWhkBIGV/ABFkBiRTgURPA0CSSHNKUVEOzwUBkGoragMmQKpcMaByBQNQIGeIaJgoakBAcoBIyfdZ0aRyiK6vmwKgVcFudMSoQmYZQId5wfuc2JmRSrXwy4wByAyjIKrGKJgYcWPPDhgJEEDVgghEc4JigGCm5hwjgcRgZUQER2gSNZZM5h1n7SwWoRcD+FZA065vdfbz+7BBgwYNGvzhQUNAN2jQoEGDXeDnX/zyP37xJ1HILKKi926uc9TFvmkZJfZDiUjETMxlKDfW1733ABjF+mVJ5BDITAHNe8/MxARpiStglueenakSUZUynpCJyPkkVU5zVokh852lef+DF86uduP1l96vBcyTs9JBkqBud8NAFhYWADBIjFHBgIjKsjSz5NgsIgCYzJu9z9AwlKUmwTKixZgcn5MVZFrYGqOqqZkRUpqEWp3OPv2pUsxDtRQYwFSq1IUSo5qm1cRElHbWvd7aH3MfsBWRtytZdIP7hQXvP3/i+B85cfxIK9+vOo+0Wn/0ROuPnjh+daP7ex9d//3rH++j18SJzg785kjJ9n41+mDgiS4cOnjh0MEvnXv05eXb//zK1X2U4m6DX3js3F9f+fa+WEBc29jYmYDeP8H1/cDdsty50NZYzPyffOTU508c9/dGlx/O8x89eeJHT5640ev/3vXrv/fRx8X+eHR8oqhnGBc7w4hpxvB11WMbMMzDTeMh4JEaDG1s8+ZBxOxeRpZBMmAAQAWwGI0QXeYee+zss89cOH/+fLdXvPrqaxffuXT941tFGVVF1UbdPKoANiIgp4E51QXEAxMQRCKmQawbCYkqNX8MEQyYnUFa55S8xGp1NEFMvyeQqxwRlX0IgIqJgkrKX1j91KmuUnW4mUUVb+YRO+wcoAYRVAAjE2QkBEREZEaXLMMAAbA2IWE0RJH0a0cRWM3KUBYqKqXEEk0RjQicY+8dOMod561Ou5V35tpZO795d1WAFOHOjdCao3/09ff3frMaNGjQoMEfYjQEdIMGDRo02B2+9OJv/+//2U+7LJeiROdy7+YWjqAWEssixqQSYuayX/SoS0gKKatfEheriKjGsgzM7BwX/b6aOvbe95hIRYmYmZJS2DlHzhEREjICERqSawXKO+dOHr52+vir73y03A3rNVtjgIaDyVs1Iw1lSYTz8/PsnCdGEBiRaxFxmg8SkaqKKjsGwGoJLQAxWzKoBkgWz8wOERE1JQ4S0zQJrXTRKbMQgIgmlVhKL1QT01CtRkdMPDg6pzGY4cA8pCF5/xDiYJb9zJlHPnf8mNvaFuAe8fBc5xceP/fanbvL+2fK8cyhgzOWvHDoEMB7+9Xug4RD/IGjR37g6JHvLN/+9Uvv7+PVm4ojrfyLZx759Uvv33tV/RlI0p7Ee2/o/mHjHrTnf+TE8T999kzH7edk51i79aWzj/7UI6d+9+q13/nw2n0yafkuYfexRhtZtDP0jZhk1Tex7FNp9wk6eIsGpx8KiacdeaGtdvv4saXzTz/11PknfeY+vnzl9TfevHb947WNjWSlkYLJOFZNxeMSekQwM1BCQkIaUsJEBgZpyE/mXJRi0wwGTA4AEIE4BaCTJTUiAqR8D0hiiqpmyX9L1BRUTaVmn0c6U7WZJOXKiBlx7jwDqqgQprVfqICECKAAmqTmZoB1MNwUFTAiIKgIALQ9I0JtnBNAIxF4h5nnPM9auc8ctXLfbvl2p9NePNDr9dU5A8NeedL6H23MuoygQYMGDRo0mEBDQDdo0KBBg12D2Zko5xmDgeeDhw61HDgG9lkpGqOYmYjGEIuyLMtQxkjEqtbvB4khhLLb66ICAseoMURhK/sBAFQ0pYhPthXsHDIAgJkRIhMzM2er3Gotdg6ePXngwunFN66sFqUogAIq0iB3fFoGbKZmKFG6vWJxsbU4vwBgMcayLJmT94YLoRQR51zqtg5nuRVvzMyIGGMIIcQYmTlNXZ1zUCdZQkKNlRqbnTOzsiyTAW6IUU2TD3RSSymJiMQYGB2ARVCJtf7pXrEVa/BJk9o1qJAx/8lHHv7xhx/KHoinwT7CIT57+NCMhZfarYfnOlc37o+X7gPBC0cOnz944Dfe++D/3buXyEz4sYdOfuPGrXsXXM8idY/6if5m6MW9CI0z5j//xGM/uHR03/uTMOfcF8+c/mMnTvy3L796vwMS9wfMYSXgAAAgAElEQVQ48Xfzm7HtU9IHDAw3NtWmk2VmXNQza+RtSlVokBjslHQPEfXw4QOf/cynn3vm2SOHDr3y2uvfefmVty6+XYYklrYsy9ixTVaHYkBE3ntVFVMQdeyc8+mXxGCE5trTvHYfQec8AJqaY4eEphJF1JSdA7MgAkCJ1EYDTMbPqqZqGs1icmNGsPQLZiDnrkXQ5gByopZzmfcoKqJEbACqaNVaLCAICBENwRSq/qpKpGSKTQginrmT5Z7NswIZeXZEC/PtuXark7tWy7dynzl0jM4h5W1x/vqdW6WpoDv3rdfvnjj8y9c/nPFGNWjQoEGDBhNoCOgGDRo0aLBrfPHFr3zlxS+6KCXgRpTlte5cK2fpMTMgIpHzGRE7j1meqVqIgsiAZAaqIjGWZYgxaoydzryqctIsiYYQJM3KzJIoKEpUU0IwA5GoRckhuBhjL3oLF86dur3ywe27/WigQ8UQDJwiEcnMJMbu+nqe5a1WpyyLGKOIJPESEZdlIaKtVp5cOMoYLWmTscovlMw6ksiInYsxioqIeOeTWFtU1azOxAQxCQ/NDCARy0ktJVEMjJAIkZlE0MDQ0nrdSnANAIi4Ryp6O/HsKF8wtmFLTEkMhdu+HW3rE81qfXLw6ML8v/3UE8fa32P2FAkXDh9q70Ze+pmlpasbH9y//jwA5My/+Pi5h+Y6X373Pd0/J5MJEOKfe+Kxv/ntl+9fEwM8gCbuBd24a4H2nHf/3rMXTs/P34/+jOJgnn2PBI2m0s1Td03PBIBTXk66cwzNO2qPChgZkSfTDo5jNLnv9mMHTpqE1P7MaR9WVlinTz/89NNPnn/6PDG9f/nyW29fvP7xDTUkR5TKESGRczyorOq0KCJ570UVVRQVAdNvEq1ixNWppRVPySEaAdB5QDKzUJRgZqqGZgDVWzOoSWdATJkHR9jnmGTOOH7u6S2BEgADEICpFkWBqmAWNAAknfbQx5oMHRIjMRMTEiBh5pzz3nnvGcwjLrRbLc+eAUEdg2dqt3w79+3c5Rl7R1UHzYzcndX1jWjC7FVvPnlq6e2GfW7QoEGDBntHQ0A3aNCgQYO94IsvfuWrf/WncpVAdDOuxRicCWhwTD7zLatYVM4y7xyTAyRm9llWuRIahjIU/X7SKKMZAIhoWRYhxBgjIkaRIpRFCKqChKYqUUIoU1q/oujm5J84/dCVq6u37nTL9b5W+Ydq20kwrKe9alr0+91u12etEMoBvZvcMMoQVdV7h4iiKqJWuWRUdUUREcmyLEmhg1ZTSqycIkFUVdUxE2LyGQEA71xaBFvPdrGw0lQRMeU8rEqaYp3QqTaJ3nkeXmOHklN248wmH0MaeeKY7avAkTINtsNPPvLwF8+cpvvmuXG/sVuF6WeOHf0n73/wffBY/OjJE57of3n7nfvXxCPzc3/i4Yf++YdX718T94AHdw/LXXpctJj/g+ee2W3qzj2jt3t+/IFjz/7+A/3yZtK53oQwPi7gJrE01tT0tlprHJDQm5IO7tTtephGJARQl2Wtln/8icfPn3/qyJHDH165+tZbb7/3/gd3VlaBiRMlW9HNVcx4ZMQ1MK0MuMxADVXVQC3ZJyciOf08IFMDUxCpQt0KgASmFiKkCDQRMIIoQFojRWAAqkZYXycFE1BJomccDyBj9b8xAIMlXzBVCRpTxkOtcipDlZ0CgQCZMEP0znnvHZNjYqLM+yz3rSxnNIeQM3lCz0AMjtAxe4fOETMjkiqoCoCRo3K9u7y6USoqYGt9o39k8cUdb06DBg0aNGiwNRoCukGDBg0a7BFO5U52eIFWg2C331/stAAgaqn9aBLNTETAkIh95s2QnW+355AIEJh97v1cKwcANZMoyddCRERU1RBRovZDqYiimuwvQggisSzKsihzZHWZ+vbzT58uEVde/iD0yyqJTzUdGyQEREAChI2NjRB1cX4+y7IqQRAiArRbSERZnptpEOlglf4QAABMzUKIIuKTR4dKls8zESIlURQixihRxDtHg6yDAMRY9SbpssA6ban8ppkQIMYYQpAYQCE5k5RlKTFWmsQxUdhWSOqv6WU20QYD7dbMBBJOebXp7bZM9FhLE9zE+NuagxgePqTPvw9IyzEQ4p99/NznTxz/bndk78iYnz9yeFeHHM7zxw8sXlxZvU9depD4kePHbvX7/+zyfdQDfuHMI9+6tXzrE+fwMMXk9z4haU5nL48Af+H8kw+MfQaAjU86AT2hFh7dNuUrHQFsnG7GicL1+0HOQBvhbxFGMhNWR01824/smBi2EOvBetshb0TwW1eFRFyR3ARHDh08e+7Mpz71qeMnlq5d/+iV119/4/W3bt+5W5RiRpaGPwQwUDMpo2o0VSQHpibRgIA4FKWpmipIBCBDgmEWBwNAo/SjAgEJCBI5DCogUrHPaTsiMCV2HCidMZsl5w0BleSVUQ9yw6VFiIAGBEAADswjOgQGIwNGZESH6JkZAREcMRMRkSf2xJ5d5l36NYIIhMBEnp13CGZo6gxRTcCYnQGGGFVBlKIoUwqERyOOVq5LNyJGhlO/++rqmeN/55XvSRP/Bg0aNGjwyUFDQDdo0KBBgz3iJ/7G//U/vvgXX4cLn+Wv98Ss18vZowhbAFVVlRgRiZhjjFEEgYp+YYCA4H2GiKBJHczee0vrWCkxw4RIBuCdAyRF0MyLaPVfjBIFiY2csMOncpfPr/bsrQ9vXLuzClUqnhHUaQlFpOz3S++dc5n3ZpbcM5DIzMqiKENZFKXLMucz51xZlmrqUl57s7IsUxJ5770SJXtFM0jm0QggEhUHU24TsZS5kJkqgbOKmqoqKoFZ8vEQNYJ0nZxzBgAaY03FzihUngm26cUDx7aCu0mC4vuPdq7gEH/p6ad2y95+0vDpI4f34D/wuWNL3x8ENAD8zOlH3rhz94O1e3Vq3goZ0Z99/NzffvX1+1T/nvBAP5Nxl/LnP3Hq4dlNye8dKYnbA2tu95hZ+7yJVt4ixDhZoQ3/IkyPl05/YGxKwXFmeesHbfMokgZa5+jQwQOPnjn93LPPHFs6WpblG2+8/d77l5dv3+n3S00ey0hpdVMKEtfrsYxRwawywUp+z2omaqrE7LwfjOtYDU2YMgYyMw2i0aqmmgogUfqp49hhVWXl4aGqKiJmZgqVJfX4GVWxVyMAD5Ah5Uy5Y05GHIjpBSMwAgMwsyNiRM/siR2iMyNTNGCiFEtHE40GKqaqYIhAhCIMYDEGQiMCIiREIjKi1vyBMkIfMRqXuHLrmZNHX/toy1vSoEGDBg0azIaGgG7QoEGDBnvHVTj1eHzb9aN2cL1UJXWoJCGZOEsU55yaqsayCKLG3X4SEbnMS4xlURCSz7K5zlyMYqrO+yzzKZ8PETtmQCJmco6JiMlYOc+ZmZAMMJotLh5udQ6u9mIR5c7qel81TBDQw2myqkq/6DvnWnmuqkl1jMkjA6DX7/d6vbzV8XnmvO/2uqrabrcdO0AIZRARAAvBA0CMEQAI0WdZkjapSjLcQEQwiDGqKiCmvgNAuioqkhb5JjrbwBxxUkqzcwqAqqmz1Yx+j5wPTpvNb9ajTVeo3SvMqpn6QNc8qrsepRC2dJreVZdmNy35LgMB/q2nnvheZ58B4LPHlvZw1KePHv21d9/7ZNN2s4IQf/Hxc3/jWy/fvybOHzr4w8eP/auPb9y/JnaDB6d9TtjVU3Kk1frZM4/cr65Mw94SJN5nbE06Txc+D9jn6QfaxJe1DSyYB8t0RgpWVOrexpRhij8AwCkU9UiXARBRzWrPq0iMeeYfOXXiySceO//kEwry4YdXXn/9zRs3l3v9UoKZGigAarKArpoiREBKzCsSEpsBIjGzIiqAgrnM+1aLql8JVafUVFQBwDvn2DFTCFFUDSHVRogiamCtvAUAGmKMZZSoapjOlUiVbKDHHj27avA0B5AD5kht9u0sRzACIwQ0IwMzSQdTTVkjpFQaaooxRkRwTI4dEcakLzcFVTAhQmaiElQlhJKqKpSIXJ77VltCLNXMO3DsdG59Cf773dzLBg0aNGjQYCoaArpBgwYNGuwdL7744v/5l3+yjBmJGmMUQYLuRg9UvePMZ2W/L1FjVEJEoqBK7BAp9ksAS+4cKnrjxo1WK3fs1jfWU7YcEVVVUMvznNmJmgIoECF6x5nnGAMAscssn8sh+/RTZ2/dWblxa/nq3Y0YtZ5folU07MCqwsqy7FGPnXPMMca1tTUics5nmSeiPMsRIcZYJvoYIIYQQ1QzEbG0JQpR8pE0AZSisNoSupoFqgIAERESIMZqmTYSkaqFICPmygiARRkJgRkVAJCcyyQGNTCbYGCmMribhWe4yYF5Qu82lRnYZr4/0e64UUbaMtGH0WXUg9dTW9jS5WP7Lk3r3ebTrAoMGPDvPkP9c2fP7NY6+ROIhcw/dfDAHg5sO37+yOGXbt7a9y59V3B6fv6FI4e/s3z7/jXxZ86eefX2nfUQ7l8Ts2H2NRn71+RuPrBfOH3KP9iUgHtIkHifsc037RY3bvPmyS/7iW92G3sQbGxPfdwsSQYMgWpHi8E2m3g5NAEZfxRSA0gEiYNGOHTgwOlHHvqBTz1/7tyZuXb+0je/+Z1XXrnx0Y1+KYieHKZlTIhUE9DVoEB1IoeKhwYkJCZWSwuUhJ3zTFUfko65UkirmYGKsjBTCEHNkFCx8tqIIqLa7/fSDwMJQUUseX9YklsbAAFIHQEYXHFDA0bIANvILXI5kJf0q0aTx5cAEJIhCgKiA0RDiMgGlPw9NMmrzcyUmQBBTdCMCVqOc88eiNWQwGfUaeetVuaYWlnW6nSo1bmxuqbK/RC9iXOt//lrr+10Qxs0aNCgQYOd0RDQDRo0aNDgnvBT//Vv/8a/83Pharv1zGpUzwDzB49oGRybd14l+UxYiNEMyHlRCyKqimCEiKIhhI1eV1S9dzHGouwDgqmlZa6hLJhY1aJhIqAdo2MQCQDILjO3YdncfL54emnxsYePrvZDf70nUxf5ghmYiBRFAYjzc3PMPDc3ZwCE5DPvES1XQBKzIOJciwhVNFHPrTxP5LIZEJF3LGpSZSaqCejaOgIBiJiZkTBG0VryWa/kTRxxPYlHMEx5iBCJKLlhmoHC5BR9Kwyn/JsFbtPKD0hhG87wt659W+uMtAW/+9zuGCa7/ECJs63wg0tHf+LUw/dYSSFyuygK0ahKiI6wxTznfce5+3ySQ+bpM0tH95w78bPHju4HAb1rPnS53//Vd97rS+yLFKKlikPKmDLiI638SKv10FznyQOLh/J8V/344w+d3ImAHnR14sVMmPf+3zz36K+8dXGnymEP12Qn2Ka3D/RzpDNfpwNZ9rndSPJL1bfv3r260b3Z6/dFSlFH2HZuzrtj7fbxduvU3Fzb7TBL+oQR0Ltknycz3u1UPmFADG8T4JzJtR8rz2gbHjMYg4Ya69Go4fgIZWkZEYBzPL/QeeTUQ08/9eS5R0/nmb9y+YN333n3yuWrZT8qoCIma2mkZK6clihVLSIREJlISg9oqmksS/5cJilkLKnFlJzQUtJAVTAVgOS/HEUMAJOJsoGZqplUnxlEQouxym1oAGaYAsymaWXQ5ivukDLiHF2G5JIlmRoYaCKwAQQsnY0aEBIjajQGBNXEtiebEBtIy5Gcw8y7uXaWu2SbLcyYZ35+vt1p5c6R967VmVvpl+Aoluo5iNAv/94rO93NBg0aNGjQYCY0BHSDBg0aNLhXhOWMTq33oXDkfd46fvSgd7kUfVNxlOZ6uLx8p+gXrbnO6vrGRn+dCJPHYhmjiChgt9fnkvI8K8qi3+8zs3cuc1lZlISIyAqkoFG1BEEQNAEAQw66qtziuY0j8/7CuYffu7Z8d70X0/LU1L9aDA0AYAYKoSxjjHmWHTh4cGlpKYQQYiREQzQAZieqRVnOzc0RU6/b6/d7IrK4uIiIIhJCIKI8z0OICQaGiKoKBnVqQ0j2kYhEFFVFVcHMCJ1zaf5rBqpqaux8colERCQzM2AGM8WYCsxEWI2yQ+N89GaqMM1IEWt77C3IxMomsyo5qtoeFLBhgU1GlnVb1dutKe6pO3bW0A1aGpFhT60JJ19s3/L98Rk4mGW/8Pi5vR17pyi+s3z7nZWVS6urK2WYenE80VK79fBc5+G5uXOLC2cWFtx+0u5WP1UGAJ9d2ov/RsKFQ4fmvd8PSe/ublNf5LU7tzextAgAl9eHPs4PzXX++EMnf+jY0oxy2icPHjiYZ3eLcuse2vjbXeNzx5a+fuPmG3fublHPaP24fzTx1NDXLk7hvdW1f33z5szFkRAZscXc8e5glh1vtw/m2YwHf/bY0owRkdtF8c8uX/nGjZulyjAguLk3ACc6nfOHDjx3+PATBxanVt6V7zoBjVNfTn0Po9HRwdsBlzxgQbdckoKborr3/pjhSPRzbGENbqp+MEgNSGtVJcI89yePLz315GPPPHP+6NGjH1698vu//y8/uHJtY6PvfEtENKqZIiHy5Ce6Ch2rxrI0AySyKAiI7EzVREHjcABL/6b/CUEFVEE1pC1mQAjMaSNoBHZAHogNwdSwNspI1s+JfQbVzdfRwADBk8vYe/ZUiZ4N0+8XtfSbIGoEMwRkYkJmRDZjMCZiYnaMRM6zcw7RiIiZO+18vtM6MN9yaCaFxOAdz3c6nXbeyh0xillQWe91i6gBogZs+e8Hu6QGDRo0aPAJQUNAN2jQoEGDe8XPf/nLv/bij+XYEoZoeLdbnDh6oN1qkRQqkQDZucw5NWjNza91u+sbXXaeiBGxLMsQo6paFDMFxKIoiqJgojSrK7p9E818poiiWhYlM3mfSwyhLIuyIJc5VobyUMedOb7wwpMn0OHFa3cBRjhoGHBBmkgHM+n1Npxnn2WqCghZuxVC6Pf7RMhEmWPTqIbeEbbaoioizOx9RswAQER5nmWZFxE1AwOqkg0mr0UVESRERFcr6USCiJqZYzazfr8wMyQkYlWJMRJikl4pkbJL/owxhNofc8dl1PUkeasS43+xJpMRAAghqbuGfO5oxZsrTRI2nF5iRJGJw06lc5iRtthRMbqZTZ6yYrua89cltqxj8kHZf/z5Jx+f20lTOQEDeGX59u9evfbOysrWS9+rjUH12kb32kb3G3ALADKiZ48c/sGjR54/cnjPauXNrQDAsXb7zML8nmthxM8sHf3atT2ntJrwCNgtJii0QVik2n5to/sPL777u1ev/aWnz5/otGep7sKhQ//y+scz9HPqvZsJv/j4uf/ipW+XlS/85i5MvLh3Dnq2hRfb4nqv+7Vr1wBgvDOb9eCwqUyFHTXIgzqfPzJT7sFv31r++29fLERGWpwuGzeAj7rdj7rd//vqR4fz/PMnjv/YQycm+vMJ8oDenn3ebIg0tlxmR9556ruazt70nBjuHLmZGAVS/HKkm5PByuRVleKglDL9mpnZ3Hz7xImjzz3z5OOPnT6wOPfhh1cuvnPp45u3e2VU4qhqhOiJEJmZiSrut26BHRMRArq2S4OfuGhmgMRIhIhoONGL1F0iUDMV1WoNlGNGJkNM+mcwQ0QATGYdqZSKWBSozTHAdPSDVn/DGwE4QDQQ0b6WnKLSKgiGBgaKBgTAQExAgN45R+SIWt7njgmhcrSu//eucqr2njK2DCKhAQF59s5578GgDKIBKG/dWV9dj9pXWP4otOfpH3z97R3vZoMGDRo0aDAjGgK6QYMGDRrsA37+xa995a//rDeOEjfKuN7tLs4vcBQwAwI09c4huTzLFND5zGctdg6RekURY0TElEFeRJKsmIhMVUV62brGmPnMAKJI3/edw8xzv98HREVg54kRrSSHSwvuwqPH+kFWNoo7vXIjio3NkUe0uAZFUVC36/O2c8zMIpJmiSEEImYmU1UzVSViYh9CAFAiq1MOamJdmZnM0lQXENPsr1psi4naxUEGIyQxM+88mIkIABIRM8UY0YwdA4CIGHFl/VEnK0wZDLe9CVuwz1PJR8RqvjtkdxEGKudqFj1x+BSydnz76IaResc4C5usZrQDU89odozRLLgdZT/12JlWju8Rzx85/PShg7s65N3V1V9759KHGxtb7B/lN6eQaKXqN2/e+ubNW4fy/AunT/3w8WN7paEnr8muvA6m4rPHlu6BgIYH4AXxcbf3t7798l/9gReOtlo7Fn5scWETAb3PD9LRVutnzjzyG++9P/MR93KJbNrT9V1Ab2ePCwMAT3RmYWHH2i6urPy9N9/S6d+i212u20Xxmx9c/p2r13769Kkff+jk4HP03bbg2KrDW7PPY8TveDRy+k3eln0GALTpXPEsz97kihkcH+A2L6jByuUKDQAIiYmOHTt67tyZJ588d+TwwaLovfvupXcvvX93Zb1fxKgggEDIiEjIRIxOIeX9tRR95Tr/YLVoKZk4qwKAY+eYidBGwpmDrhJx7bxVEdBMjDSe+DfJnEVMbDC4VsLnioAe/aBVww+COSBvRAoCWqIxIpiaKiMQpoUCgICO0CM5xMx7z+SJWpnPveNKoo3p3AhTpkRmRiJgUJBy0ENVLUMZIxiAAEopyxvdArAX5NCB/M5KsfN9bNCgQYMGDWZGQ0A3aNCgQYP9wRf/09/86l/7ub5FC/2PlpdX1rrcX5vv5J7JNCXVI5/lwA6dU0CMMemD0vTP5zkRJZ8KQOTkQRFiPHDARAhAVaNIjDE5G66truWtFjHGGGMIZVFqqZ78Yw8dFYMQypffu1Xe7QKCjMztAGp61ExEil5vhe7Ozc1lWbaxsZHneavVWl1dRcSFhQUAiDGura232u1Wu5O46TKUzIyAqhpjBDDvszR5LsvCDJi50+kgYhlDmoSKCFICgJmJCUREzLKs6g0ioiKi9x6RYgxKqiQA4JwzlShRAUC2MeOYnPQbjGxAHC6zHvln9B1CNUXGkfn2eNFBS9VcHSpaYArXMCJArv6xmtIeKt1qqXI9+YdKO1ZXWJMNNiZSHbX2GCwqr88SajPuqps2dgoDlmFzh6vaB67c+wpC/FOPnp69vJr95geXf/vKlQkOBgB2ckWYci/uFMX/evHd/+/jG3/h/JOHd2lwXHORY5r4z9yD/0bCowvzxzvtj7u93R+6WT+725s1dqCNX1VM1BQgAPRFfuWti//RC8/tyKU9Mj+3uYm6qql93gv+jYcf+tc3b14ZcQuZ9kiMbtnbYzyhfd6Xz8LUh3b0odpzaMQA4GSnPYvbzP/27nu6naW+AWwn3e3F+I8vvf+tm8t/8cJTB7MMZuLH9x3bnOY2vPPolnHeGQY2TJstkiZK7tiB+w4D05q3dZlfXJx//LGzLzx34fQjp9ZWV9+99P5rr7/50ce3RKDbLUpRl3kmBjKzlMHPsDJGBgSkZApdhYopnRsBAhJYLXw2UJEoY1J3RCSSpJAmIkYCgBijxoFpuQFWSQxVk/+WggGoJB9nMBiwz2mEGjhBM4AHypCcAYCImYIRAAEQO8/smRmRAR2CQ/REeZZlzJ6IwdIyssqFg4mZHA3SEiISGECAiAyIGEVUbX1jlZCAXT9Cn0jYRbDFOF9Q+dV33nlQ97ZBgwYNGvyhQENAN2jQoEGDfUM0ZYJQFkLW74c2Um+lJ8V66Hfn2nPO+RjE2JH3ebvDjgFRoiBRnufMlByWk30h1TbKaDpQRjEjO59SCDGhmjExgIlIWRT9EItokTLnjs+1O2V4VWK53I2lQaynejbknRDMJEq/1yMiAEgi6I2NjaSDXl1dhZqsLMsyigJAcl9UreZ4qqqq/X5BzIRYzTbNRISIiqKoJFJmCIBEjsnUyhCIkJCwNpklrOl1ETNQkSSeMjVTS+qlGGOp5dCJeSsaxaZQDxP6rfTPFCIBcVQkm9RY2wiTsaZ0p3RhrPVkjA2ICDZOatjQ7HNAO4/q7GoRNsImrq0ysB5trNJ04xSSZfw0BzsnyejBnh3E5rvD544tnex0Ziwczf7eG2++vHx7C65nYqONb99SyHlpde2/+c4r/+Fzz87YjZHKxyTwZxcXlto7i4J3xOeOLX3l/cu7PMhGujSQ2e+WEcNNL2C0tlFK+9Lq2vtra2d3UtceGVNJ26aqJlrc46NFiH/uicf/1rdf3qTh3fITes/YFNLaSw3bH3gv7HOFWR7I5X5RLybY6i7MFCF4b23tb37r5X//uQsnO50HroDeSY+8VUkYC9RVG0YGkhQhxInyA9iWb6ZsmDkkZBN9rMebqppBLLAyzDBABUAiBCBkPHjo4BOPPfr442ePLh1ZXV+7+O6lV1557dbynW63jBFiTGN1VDJENTDFiBjM0Oo4qyDSeFSyztZnZiZERAwAqqo6TkBDFTSuFzZhKlaPJlWINv1WGOikAVJWTasU0GCDiz74QDNgC6mFlCE5QAJCBCJ0jI7IEScjEQIkBAZIL4xIkjmJGZkFM1IjVEKoTMFEEICZHCORAQUiJYL004II0RF32rreTykn+oBI/Xndh+/5Bg0aNGjQYBQNAd2gQYMGDfYNX3zxK7/14hdi9ODUQjQ1EQ0bG+X6XTiEeZZtbHQFEJ3PWl3nmRDKMhBRkgybmag45mSajACEyAxMaaLHRI7ZMTMhZVmWVqM6x4ggEvpF2S+DGCwuzJ9YOnZ7ZSXE+NaVu3f7oRdVARRG2GcEAFBTLYs+ESItLMyLaPKAVtVutwsARJRlWVlK1MIxp04WZQlm3jkAkMqyAx27RKBHERUBxBACjM9vHbOpFmVI81YiSvLeRLcbQCGJ09Y0MU7TSyIkx2ZAFCuFOMA0CqHamnh2rLMuTuVTplIsBkBE9Sx64NCxNVLypc2ba21yzRwAgBGS1frqREbXbyeZlCrh4SjLhnX6JhiZrCPCuMvGkJwfV7VO9HF8pfceJLS7xo+ePDFjSQP45Tfeenn59vbFRjo92v8d6LO7Rfl3X3+zkBmNa21qhbOkH27E8nwAACAASURBVHxvde3s4g6k7WeXln7z/cu7ufT39zbhmBv0QLwM37q1vCMB3WLuONeNEcY/M7bfj9fp+fkff/ih3/nw6sT2rYntXTU+GszY96s9Su9ulmzvFjYinbZ5v3OuwtVyIkvk6FfP6Cdo5/6slOXffuX1v/yp57oP1AP63tjnidc2iLnUO+pvy+0vwE42UIOY4o6lNj1hY88F2sjiF7TK/JjS+EDUmescP3H8wvknH374pPPu0qVLr7/19hsX35WAZWllGQEIDCRGQAFUpNoBA2jUVArrD75Zoo+tWi1kCnWE2Ewn45GjS3KQJk94EAEdyu2tGp2GthvjX9ophSGAQ2yxGxDQDEgIzpFz5JkIKaVtqOK5AGCgYKoaVREUAcmAwLAKDye6XdGMCL13TlMixoikjmE+MdCOXWeuVI2Exq4syST2cvgHL720841s0KBBgwYNdoOGgG7QoEGDBvuJn3nxn/76X/kzsuHacyqsnbzVXpyX7jyBgUgrd0XUILHod0OBgBBCaWrd9dWBD0NyZBSRNGViBiIiZqxEP+ic9y6tQyWoPJTZeyYi78gZ5I47vvUTf+yHjh5/mP+fb7z94fJHdzbG6Ic0FUzzRtXQ74OZd+x8lmXZ2tqaSPTeA4CIrK6uARESF2reuyzLACDGWPZ6gARESCDRSiuJ0npcFFVTjWVw3jnHRJxyGKoqErXbrURkxxhNzUw1mTqmnEhKyRSbERlRJCbCGgDYOYvRVAbUan0yAwwmnlV+QJuYGw8p6yk8woB7UJ3CD9SF6qk1oiWJ+qZODAqMblCremRgaENjTRwwf1jVX3EcQ0vQUUdqGFAllnTlA5H2iK55QGRvOmcbMNwjF2ET3WYjp3nPeHRhfvaUfV+9fPk7y7fqXsE0jmzTm0noNqrSj7rd2ToyQZFUfSCkH1w6uv2RV9Y3fvfatV9afGr7Ykda+eMHFi+urM7cnylbdi9/HlQ1IXc1m9TmV2d9fTafkJy5G0N95LBX40GgfXicfvb0I9++tbzc749Wu+k6zESkbjpkavfusc/Tb1z94h61z9WLnHjHY1puUGb7MxqltrfESln+8htv709qzx2wFe88/f0m9henJYcd/B15UBHQRujnkYOGwl6Awaqd7bAjR40zPFWWPpNVrgKsvs8NwMjRI6dOPvXEY2cefYQdX/vo+h+89M3LH3zY7RUSTARNsf5+AAQgIAJSUFW1SdNqs+QubbUwOT1LZmm9U/V66kBQjT31xRnjnXXygpjWPRp9em30Q4AAjjDzLiPOgFiNDAAM1SxICCEx8gZqZqPmUsgpQmsMxIm2JmBCImZCR5RnWSvPWu3MMTEBO3OM3lGnlTFREAlEG92iNIpRbt7ud9r+n37nzR1vUYMGDRo0aLBbNAR0gwYNGjTYZ0jhfFaqkmP0TAtzc+QBNEoMZcnz5IxclDSDMolRVQYLVRFRRWKMptGAzKgoBMzIsWmaLBJR4maTDIgI0XnOWzkzVqn1yKNrdVoHzp44/CMvPNUvX7+zuiE1bTughLBW6apqLMtut9tqaZZlC/PzROS9BwRVLYqyFkMhMznn2hJjiBICMhMREabEifWCVkoEtHUs7a+X90KM0cxqN2gQiTGKqlJKeKiaUhiyczWRjJhcRsCS3SQSSsQYBWwwxcXReex2pM7oDtvEQABUfpjjkuGaAyYYTHphhOYYOjIP3uHmnE3DIuOEXLWrIsyr7iT59qBztXkHTMqih923SiKNI22MlbEB2TzCBU7SWJPYJxeOz584PmPJDzc2vnr5CgDsnpjbXH7P7B5sQyBdOHRo3vvtD355efnV23eCqt+Jq/rcsaXZCOiJEMuoUHcPwJEXEw8FwFjoxABwk3J2OjLepjObW9w7MuZffPzc33n1tW1L7QvfjfW/9/5B2Meqtq5+WxzJc4cYp3+o93KD3ltbm7HkPWBG9nkYgBvlkIdlxr+lJ7TPA0xGKwc1jIX2qrFs215vTzBvkR12fMxIzSKktAlpZARkXDwwf/zE8WcuPHnu7JlOZ+7SpffeeOPNDz64endlLQRRAQMC5tGrYAhG1YhKTNVymmrAwuSahQgIDAZIBIigWvPtlH4lEGEy16p+NlTXNamREQGRKiLbVFXFtOaXU8pjQ4DaecMSA28T503VyiwU1VKVzdAMKwNoQzO0xMdXqSCIABGRzGEy0iCP7Il8cn8mRADH7Jlbmc9zn+WZY2QGZGNGZiJAAwpiK/1+oVCq9IDn53l9PWx7gxs0aNCgQYM9oiGgGzRo0KDBPuPn/7sv/x//yZ9iFoZoQI5hrtMmFFPpF0Wrs5C154pSRERN0nwtxhhjVFVCKsuy1++VZYmEPsu7G90QBARjFBUjdqYaY980KT2JGJ3nrJ8ZSJr4mSGQay8emmsd+KHnn7r84Y33rlwv+qpasbZWTcERUuI9NFXtdXumRkjHjx/vdDqQJq5mqaMG6JwzMFUFqCyaKz9GsH6/X5RlnuWJWQ6hNDPvvaqJSFkWzJx53+v1Qoiq6rwnIkQIIYoIEcQYy7JIol7nKhEWAhCzN1DT5AXJjkMZVPu1FwcO6bNaElrPa0f8McaYiokNOCgOQ7q5FnNhRcghspngNFoBK7qh2lcR7gMfj9E/I41X8mcYkNZo1ZwfEGvi0rCa3cNQBW024EkGf2r12eBKVJWPEN841LQO6fHNbPVQHbs/TBkCPHv40IyFv/zuuzrJzeBon0Y2bo9Rbe9usZUSFgDws8d2kD8DwHeWb5cir9+588KRI9uX/PTRo7/27ntBddtSmzsz8szfK3DotjHC2Y5y0Dt1r4JWpNKOoux9IGEvHDr0uWPHvn7j5rYt7qqV7Tt/j33e5nne7YM6NRSBQXe2wsiYzx868NrtOzPfoP16xvaGyW/q4d/R4MKom8QYTTzcPChpNjLuTWsLp7guYf1/XWLwpbr9N+SWV64eGnaisBEAAQkZDEwDEJAjl9Hxk0ufeuHpC+fPHzxwsLfRe+31N7/+jW8WZUiDNCAhMbIbzSdpAEoAZkBGzrEjIlI1AGCmGGIIgZiICDGtvwJETEt2mJkQAdExq2pRltW6qWpgQkzHABATAKholCgxaoymViXFTesrRtjnMYa+Dh8TIBmpWiECURgM0RCAq/+Rqn8REYiAmZiBGPLMZ84xcYu5xS53npmIEFSZKHPsHTtHqTwSKCoioElRinG+sl6sWyzI9REYTHL+2qvvbnt7GjRo0KBBgz2iIaAbNGjQoMH+4+f+y3/yW//5FwJlDnSjXxw5dlQlxGJ9zjvnc2KX51yUQQphdo6R2SOWZppned6SVqstIsTsM9/t9MsyAECIIlEAERRVLcagqhVdixBiCDGIRFNFJCLtr65YrxReP3Ps0KfOP/b1Nz642ysCgNbsqpkCICIlhRKIlEWBiN1ut3JirlMTAVJiYWsNsgAAMyc5MwComqnFGLmCq2hPBCLyPmNmdjy/sKCiIsJ18h8REVFEFIkhBEJK/hApM5CZqaiqiorEEEMoyxLMwPIQUGIc+jWnMwIYcsRJp1U7X45sBJg2/Z9CCCQ9edWEprn0WOkBy1ArjBFQzRCRkGBEZYxQU3qb1MkDQsWG96VipmhgwVmVqHo1uvq4olQmZXk4bKqmXWrBuw3KjwgHYfzE9g1nFhYOZDsb1ALAxZWVdyo58LRbUZ3GkNYf8fjeVHak2C5JtCH7jNUFGlaVMT9/+PD2x9/q969ubADYt28t70hAtx0/f+TwSzdvbd2ZyS0D5eK+8IOjXs+j9Q7eGsBitoPiO6EQmc0PZH9ozS+dO/v6ndvrQeo6t8JMbSHC0IFkCqY+ErNjm+d5dO+MYZXBBRx+t3TDTF7MP3369Gu3727bq8mnYLaO3Q+MhhUBYLBkxcaS941851n1nTB6i0bDk5u9mSfPq6oYR3eNlxkdS7a7KtvsGy5u2VxoWD0CABqgASGCcxk5aM9lD5068ewzT73w7IX5ufmbN2/+wde/efnyNUSXt7xV9hSYLDcGOQMMKqdnBESDNIITUQokExGTc84TUbp6oooA3rsUPI4hIhEzCxoYOvYGZmApSUNNVgPWWQoQDZGIGcA0RBUxFTCFFCOp2efRc2diMANTj+jAIIgjZO8ZkBEIgazioAmQEImA0AjNeSZGIsi880xMlHFKVEiOiJCAyDE65izzTKgqZRkNlD2KaVRD8qLSFxFyRUQ0lQy/8tLb29zaBg0aNGjQ4F7QENANGjRo0OC+QIl7OJ/Bek/L26trc3Md5IzJkMgAidl5MEPnODGD3mdq5p1T1Zi1KIl/wIi8iKja0KhDzQxERJNpI4KqloFDYInBzAiQiNUgSqlip5cOlIof37xjN+/e6YeB8rYy/ahX05qZSCyK/urqagglpZR/lrwxQQESO4xEIgIAjhkJ08ak4B6opQAABpwoIhOlhITMjICiQiLJu0NVVS3Nh0UVCQFAE+2dCOghTCxpuJG9S2SwiVjFCxtMEgzjtNH4vhGXjXE5MQwICBtok9Nce5i6EcYIChylOcZqHpRL7P24NG9TN8fXbW8iRwZnM6qh3FzNsMxIvQNKpfKhBsPxy7VZzTeak+4e8MzhgzOW/BcffbRTEdtei4pj5JCNlJ+RQZta87DWTx85kvEOZrvfubWcXry8vBzN3E4uuZ89dnRrAhruqwq1plO3axsADuf5jlUF1fWw86L1HVucHQvef+nsub//9sV9qW0WfFdY2BlxuyhmKfbowsLPP37uV9+5tG2pAQtr9/Xx22/YQME8Qm9aZe08yfVvgQlif/Mhw6x629aCs1y30SGppsgBhpbKAICoBgjAiK2WP3L44FOPnzt35vTBxcUbN26+c/Hdt966uLLW1Uo9PK4Bh7Ha0qicYrqgJvUaHR0YWlidiVDVEKq4b5QYIxGCmUapjJa1yldY8c5Y5wVErI7XtBJLTaJJBNPq/4p2H+H5AQCAABiRgNrEObJTcESOOWUgJEx5BYEx/bBBIkQ0IvPeMSESek7hbCAiIFJAAQREIlSAoIoiKBDKUjQiQQszBVRkJe72y+A4hhh6SB5/65WGfW7QoEGDBvcRDQHdoEGDBg3uC7744lf+p7/2l16Xp37cvnU1rh8qw+HFRdCiMjQkcD7P8jbWSiIiMoMQShFx3rz3IYT19XXvfeYzUyBGrBhbVVVmBgRVKYpCRIjmTFWjVLnpDMoQi1J7weYXFrKsdf360TKGtY/uRtOU6bDqaG0gDAagJiHcvXO7KNqLi4tFKGOMABSiRNXMZ2YWYkzHqgokBTVxIsW9cyJS9Gs2BAkRmbndbkmUsiwrA8qqWQAwVQMDn7n0hpkRQFRVNDliDzoJaEioImjgHLN3QBjLUkVqx4mKbBi6G6cpPRFWgrAhQYnVCmUbSLcG1EIlF0vUPkJlTE2sSgAwwrDXqmcdoyTqGMHAuGAHHa6NMMWmZmCDJkzVYCRLYV1sWi1TGjGzwZLqRC8YTqr7avp+pJIB5zom2d4jGX12tvSDvRhfXr4zfgI2qkXcZGE9Sdbj6H0HGFF2z6iDHtBto+kXx479zLGlHU/k28u3AQABC9E379zd0X4kmUpPY28HTQ8oJIChvv9emcHN8YVhcs1BAwgAcP7gziGEm/3+6IdgagLLfYpoDPFDx4/9wY2bb929O3KvYfSWzZ4iz3bo/OhHcLdXfoQMHenV2Ae62r1NzXXQcIzBx0FV12dNrQk/evLkiXbn1969dL3bnbxckx/yyZ4/WGwK9W0VHtr0rTet0OZP82iNOLlhy687G8k9sBW2JaAHy1yGHR0+p4PFLkQIgMklw8BApdOZf/jE0tNPnltaOrK+tv6tb3779Tcv3l1ZDdGiQowBDbASMVt9YHUmiMCQ8vShqo6OOFhvYaJEHqeNaWBVNTBTorTYKO0yUR1kzcWae04DlimYmgqoJm4bTEco9TH6fvgcqzBRi3mesxayN2BOuY0ri2lKV41soIBGQiJMKQUJsU7IDIIEgKJAAITmgUA1hsBFUNWyLBgxz5z3zJmPphtlCMglaBeCyziWOyfzbNCgQYMGDe4FDQHdoEGDBg3uFz60h57zH/h2Fta7tzdiUQbSsuj1QGFx4QB7ZwbOe8eOmQCACLM8S1OpoiwBoNOZy3xGgDEKMQJBsoo2UyI0M1Ew8zGiijIzOgeqEqNEaeWZd8BFpJZjn//wC+dL4Dvd3q2N0IsplTyMEnfJ+wLMVCXGUBSFy5z3PkQB+v/Ze9MgSZLsPOx773lEZGZV9TF9TU/PTHfP9OzsHDvX7gDEihQpYQUYlrZrhCisBMp00HSYTCb9oCSQMPLPyGSAjEZJlImmgzJKRpkBgrRLCQSWwgJjoLCEsMAC2GNmdnbu7rl6+pjp7uqurqrMjHB/Tz/cIzIyK6sq+5rZH/F1W1VmpIe7h7tneMXnn3+PWM0JA+ScRAmUmVhtExktiplYOBBInItPtswsIlnmggssJOLMzHuPhu1zIOIscwCCKkcS1jw7jmRpFHxrUMDMVJwTZiFiZpiNmKuyrKqq0UG3LAXqZ101g04TAjSJN1WHFmztCqYpKjPla5EdMPAUKWuJNUieG3U1eBKArn78nseHNfxv2sYs1LaZJpZIsFgdG7HFJrcyaeiV+bRbE29xwqK1OehJNSNvMksc3jT5bADuW16IgH796lU/x8d2QqPMHNwx2a1Q5tuWuJJnu1Kxa2X59tpak8OLly/tSkAL0ecOHfzmuRn1d2spANRmz+pPb75XUhZbLzJxSpNvkBly5scWsPA+s7Y2YcrncoDbHLxF/PypB3/pe9+vNMztMpvbmbugbe1L8w7eQJ778nzHHQCJUiYQEzmiXGTg3Jm16+9cX99S3KzBTrtW16vqyni8iFYdwKf27f2bzzz18pUr37pw8dXVq6HePrLjVX08HDRtebn1SHpD2yabuRDClNZ4a1Zz3m+LOT4eN4i2hrpmiLe2vDbG68S9XnHwwIFHHzn12CMP7V1ZOXf23CuvvHb6zDuXLq2WpQVDiCpmojhlaj1ltb7TpKRMTBSn9wDTuDxMzX4jGFQteLDE6H7RLoOF4t8EUK8AkWxZrElxGdPVpT8q6rXg5kppawRdRFH2wEnPZT12fUhmxEFJQTDETUftjRNkjdTbzMZlBTMii38RAGACEUwDMTmm3GVMRGb9XuGyDDAnUmS5y3tuMBhubHizseoYdHXo9/XxjbfevqXO7dChQ4cOHXZDR0B36NChQ4c7heeee+4P/5ufG48ruHw0HA5Ho4IwXF8fb26MR8Mszw2RoWVhZ1DneGlpWZwA5EMQdr2igIKJvfdRAR1CMChg0aG5ic5nAczsRExDfPAr8sKMiEvOqHD5o4Nj10bj1c3NH7x9/qNrw1Kjs3N8uGu2KifjC+/9eDwSt+RyMYCFLTGtBHCK/1dLtJxztQDKADggy7Jo68zMzBJ5UxFhETOlkIISAVFAHQPsYRIUMXpAc1QzqYXATFr73xqg8TmUiVmYhUWjDrpNxLZg0Cn/jHhoHu9AQOMbPTkCm9DU059OlGw28XI2YmoxJFwT/BPmeqrIpG2NSq+GAbbWh4lGoJb8uv1xwzOgzbUkH45EchBomlqjViaJIIiBouaJY2+S7TzQK5azhRyE37h27WYKWBS3gTv73KFDvBv39NKVK+0R+OLlyz9/6tSuZz17+NAWAnoaU+1/B3jclO2civ7M8fsGbvc/lV9fXbD7ZjWot4hD/d4Xj9/3G2+/c2vZbC93vTWi/5H9+x/Zv2gEzgb/x1tnpglobLfo0sZrq1c/f/eRBYtgoicOHHjiwIFxCG9dW3vj2rUPNtbPbQyvlePthc93moOefzee1wEtT6F0gLacYpPjM+7eU5x2nVVt4r9bHXkBBTR2aajtFn+mTrQ4Fff7gwMH9546dfLhhx88duzo6pUrb7xx+rvfe/H6+mZZBXCmoLS5hdk0rSBb0HoutZq1VYOA2DRAg2kAM8BWTzdqBlWopnXI5kqjM5RFOXP0fua2aDv95WA1tz6hnds8u83cwuL5QpQzD7Js4LKCJQvEmmZYU5ikP0kURtHcmsCKUE+LwXszJZiIix7WLGCCITgmFlY2EZdl0iuyzDnNRFiyvMgHS2O1kUJZKuPf/N7LD9994FtvnVugZzt06NChQ4dbQkdAd+jQoUOHO4jP/ydf+91f/tlyYwTyEGKm5X37oNXG5lrhi15/+drVa2VZMhFxYpDjI58SMYuTLMbXgZk4ERHnHDgqXZmFnJPofyicfBC9ssuKXl8yyVTNiANAVK303Wcff2DvoQPDr//T0XC4OgIzG1GIwiagITrNzFd+aCMFCu/zPM9EQDQej72vvEUtFcEo6JQ2MIQQt/H6EMxs4tFBHCMaJQkvU7SYVFWCwZTMQAIRFgZgqnmWucwxccyNCQDUqBqXplY/HhuMiMCSpT3HtXCMZx555wQAtBm5KyOpqNqP0YRIHEdilgBiIjUz1dgFxNwQxhavVgSAESyZd5BpZBMQheMxFTGnFzXH3Gjj0sZjg6XN1BqdNACoKdSakIfMUQ/GUfLW2IloErg3lUpP9PGKagGZmSZuxibJor56euP7DYtXU7lH+v0FT3hvlnFrMCGg2qR5UzWacqWYPmGSw6IVbrSlmHpDAJ49dHjXXF66fCWeF+uwUYU3rl3bVTd9YmX5yKB/cXM4XWdL5M5sxWpN/PSRBTEh7mbbsVnpmFi8PLR3708eO7ZrnkPvX75yBc2XbKfFixnicCesjsf7F5D0fuHYse98eOmDjQ0AzTJQvQyweGm2ZXSl4/Na/s6Cp3YlzGFg6xCirQOwly5fXpyAblCIPHbX/kbkvun9xc3hh8PhheHw3MbGe+vra2U1tw63H9t0VHtjyiTVjM/+1LCKk2P77fRImCKuiYhr9nmxGwXxrkkszk3bgaeqWp8DEFicqsGUYURGhHvuOfjwww888cTjg8HypStXv/WtPz5z+p0rq+vBq5qBSqRYEQiKJlitqdUy5FhEMIOJkokFb4lojkut6XI0eACIU4maUtrKE0MWGzE4r6s8YfhtanoIaZKJoSnS2uzUOG0GdLx/ZczLzi2JK4idKiz6UZtxirygpiGE6OZBaowm2zhjGgNCKHLNMufEZc7lmeQZ9TLXy0SYiizrFb0iy5hFvQJMrtgc++u+9MLjSlevrD917OgLH+wagaBDhw4dOnS4DegI6A4dOnTocGfxhb/56//Pf/ZTPM5sX6jAfeEDR476jTUEBdAvitw5gGLIPR+CafSLEFWtrKrK0tSinQUzO+eitIk5hgQEACbKnAjHGEFwzuV54UTMEFQBgjjLykG+dN+Bpac+dd947F86/WFlGoy4eUy0xOdFgjN4Px6PI2G6tLzU7/eXlwbBNNTPt0SswcwQa4L05Gu1khaqyZ2ZWWIwwdQiRBpCMnrWoBrUByMCMchMLRLZ3nsi9j744Ln2ySZmwBJrYEZMceexwDRAERD1YDe+ozzJrqbYKzPM0g1ReF4nmrOteFLChOGOjQNirgMNJtVz8zOyX1OW13V4Q4tdnTIhq7eBJ6LYWqqzdDz+mFA3qgZKI2zClk+us1astaTXkwa6GfY5YRECMZ5wblsT2ya3+fSQzSa7RczmE98f7veP72ZmPQrh9atXZw6+cOnyIh7KP3b40NffeW/LYap/Nn3S1Gorh7UwtjTVHLIOePyuu/6dTz8sCxgO/PGHH1aNLHQn9vnG8L1Ll+9dWnp4396dkzHRX3no1H/1wotNQTddYlp/m81gKuM7zsNGl/mpchfCy1euXB6NDvR6t1L0wLmTe1ZO7llpjqyOx29dW3vz2rUfrl69Oi5vJfNdMMfdIt3fmjsR5psrt9dpkG6jcxrPaqoaU2x1uh8vuLKwwNetllRv+ym1ljNQ32ApfQ+FTX0gpuXlwaGDdz3xmU8/+ODxXpGfPfv+W6fffef9D66tD4myLGcQjCLXa1NZATAwC4HSdBwnSWJjNhHEKBGc9hgln2cAgNYroLWe2khka9QBa2b6JJ02mGlQa9+itpsYDTAIkBEVLIU4Cqa+8qamagYzaFRdE5mpmgkRm5EqE4RZnMRQhMzimBxzkbsscyKSOc4yzh31MimcRBeOPMtFGEYGNnEV8eZoXBmNS7sWqL/Ux8buvdqhQ4cOHTrcFnQEdIcOHTp0uOOgsdiSkYh6CkL7l5d4MKg2N6vKL/WXmgA+la+G41HycAAboGq+rHwIIQTvPQEVi9XBgmAWVL2vACsyB6iZgThzWV4UXENY2DlzGffLwvUePXn3tevD9z+4crXUUVAGhcmzfiI9I73rqyqSkv1BL89dr+ixiMJ8FdSM2SWlFyXRWduIA0CMbmQwiXWO9K6aqtY/TFXjpUV6WlVD8N57H4I2emFQpLmdE2G2LYYSAIgQmAyEEJKOCqgfyycvd0BtMDIrLZzpyaQ1TufA1JoIh6286jrNEIVE0Spao/p45ixKtpwx9BMITByrUNt1wpTNNKqnYwNORRFMRddHGqWzGU0CqTXJrTFCmQ3b2Mppl1abj3TWggT0RlWNw8QAei791tYx2mwy2+HERbp/5xIBe/bwwZ0uAADwwyurPinKJ/LkFy9f+VdPPbgra/XsoUP/5J33trZ13WUTymrr2sn2XNccTOUyf9DiQNH78onjnz20+yUDqFSff/8Daxm3UGv4z6qh50mkd8D//uabf+uzz+S8i+b0xMryXzh2z+99cG46VODiICKasX6m2RvMxweelvnODACq7YtmLtaA58+e/flTp25vZfYXxbOHDz17+JABb69d/85Hl/744oejsNWu/XagvfViQjpP1vDiyovNytB3WDNASwU8w6PWU8ONr+AshJ1XblrS59axyCd7Rijy4tCh/Y9++lOPP/bIXXftPXv2g9dfe+Oll18fVwZIXuQiDCIjDRaCzbGTt1J8SgAAIABJREFUcpIB5IOHgYgkcwBUVc0RwMySCGhWVVVjTlYekbBmTv5azMw8m7mZhZAm8TQNBTUNRlp3zZZOmZ5WGciAnNkRW+V9CKTRRMsMZASjJOgmgESEwYbMSe4kL7JMxInkuXMijjnPMifCQuLICTJGJpwJ58wiTkTSlREp8/pwWAGjEMK4WhLZkOyb77y6UJ926NChQ4cOt4yOgO7QoUOHDnccX/x73/it537GFOQsEG+Ufu9gz/7+ysrS8vr16+W4BJFaqLzPxiN27DKnIYzH4+FwtDwYMElVxZ2zRkTe+6qsLGiUIVGvD8AseO9D8GYWqmpYeWKa7EcmMhbPVzznwsWxff0nHzz82tnVC1eHJSEYRVaVAVC9f5YAM/VWQq+u6nC4meeFyzKOYiIDNNIhFGp1NoAJOQ4LQRsSvCGg037pqN4mJiIRBhzFuILxIVlDfBjWJGc2S3R0dL9IRSRXClUNgXMXQhjTSCvSEDREUj0+wyYPjTYa2q7RCTO7JKyeIo3n8AhEqG0sWtxIjYa4mqHjYQaFUs0QG2w2dppBCUTxMgEyTlQ7CRNHHw01VSBMeDxLO/Itss01U9Mo0YnA9aIFGNRcnoE48elzxJ+3g33bm+eLJFsrp5SVc0tuKHKrFeM2W2faVnS3G7Zqglu6RGAx/40XL19u+OK6VrRWlqevrZ3au2fncw/0igf37nnr2tqkBrNcbRqLNj3aUqiwxVCIHF9evlaW16uqcUwHwER7suzwoH//8vKTB+46uWfP4qTcb79/dq0qaasnyBRJaM0mgBuBXRqNv/7Ou3/5gZO7Jv3S8ftfunTp8ni8ZS1hoSJ3cuX92EFp+Nh0z9a66MQ2z44NAH944cM/d/TovUtLd6RWwAN7Vh7Ys/LlE/f/0YUPf+fs2etldScK2lLsNGzLat92Z2w9tblTTG6BrfvzYljo27ZzltNU7ETUbaahJNLM8cnj9zz+2KPPfvZpA86dvfDCCz88d/4SUZY5IjCDzUyhRhARAnuvMxfSvLF6GXQyfcaiiSy5YBGAsvKAMXFQBYyZVS2+iPbKsxeRJr+4YSoACmhtFR03Bk3MstsrsVq/ZTP4oMqiRkYwAZRgDHLOiYtbnYiZMyEhsFkmlDnOYiBiJicQViE4eIGyUcbOOSdMzMxERqJGplZWwasF43E5HHrbDNgYh1zYhfD8K68s0KMdOnTo0KHD7UFHQHfo0KFDh48DX3zuG7/13M+QcGU0qqwfdHnlrryX9X3InAOxDz4LPisKlzmXOVioynI8HjtxMPY+TAjoyldlabUAlohUw2g0DC7EmIQ+hLKqoqZJQ1DVSEKrH3stpcCRld7Tn7qvrKzy4cPNyiPFIqqJjQlnahaCt+FQS1/lWZnlucscs8DI1JgEQOUDi0jaq2uqFgmpaBsiIkkKbY2kCXH/LEkkkeOWXxYRACIcND7xWgghUtbBB2sqGO2kmWtPiUhSawieiSoufVl6g1moRc2L6txaD+21CLH5bMJsRfFoIx3WlshuCkRsMMTGJyIia7TJIHC94bnV1jqhUaPeOYnSiBJxXBPQjcqMiBpGalJda/1uyyQpBkJs9NFm0xrbZNOByYGbwOS0QmSREzb9jQkqb0GavV1+2+VmAJ1cWTnU38XZwKu+fGW1fVqDFy5f3pWABvDjhw+1Ceg7QYAe7PX++tNPxtdq5s3UjIl2lRhvh/fX159//yzq2k6+Pphp0ZtXmf7eB+eeOXiwbQoxF4XIV049+D/+8JWbXoT40YFs31o7X5ua/W+vv/ELTz150x26CHoi/8Kxo5+/+/A33jv7Tz84p7dzpM7In7d5ixk6dLq9iLYcbryH2ym3Vvs2aaEXbo/EPgNxFZHIQLp37/LdRw498dgjDz5wot8r3jrz7htvnnn33Q+urQ99gMUJIq08q5LG+3ecYduZe/Mg0hSrgHzlQTCzoAqzEIIGJaKgFqvhg4KMKQmfiTlSzCRp186cC410toXakkNTYIbJ/7RsRq3WZyAjzon7xAVLRiLCKfZCbAeYcyJOiFBTycZkQpYxOWHnxAkLkTAJgQnCJqREZBqCt7hCWyXfKSaWUo3zfiDa8FVl8CWCk9KH3+zY5w4dOnTo8PGiI6A7dOjQocPHhC8+941v/PIXXTb0m3uuj8b9ssygmeOe6xHRuCRR7rssOk04BhPMrBxXVeVDUFMQIMzB+6qqYvi1KGIqx2MwotmFOFeW483NTREx1ejjTMwuzzPvufRey4PLe44eOXp9fbgxGl4drfmgRk0Avy1apyiFgicSYo72IExE0dOYiII2DDK1gtiFEJJ+KjHFiiSRttaG6EYRnHTNNUsbye+kdFZTZs5cFsXU3sd4hlBNEq3xeMhMmWRjorEBaiFYqC1CFukdteQB3U7f2gHeqNSUWepqq2ogcdNKRUrnMJGamsbtziSsQWMjEBML25RsjVr0dnrgT40WTTGpaSdDsodOqtIm9mB7k3mbRVYNVPuAWoqRVbPX03ptmE2E21uErAtgKnG2Ze/2XHjVeYe3o8DnC/1uli9vs89NiVMLA88ePrRrLq9dvToOvpXDRA38wqXLf/mBk7s2xNMHD3719NvVbFNYSwtNLZq3/vJs4XoXBBPlC/g774CNyv+D1163ORLSHb5xU5VfAGbAr7755i8+/ZTbjVR9/K67Pnfo0Hc++mjhzNu12q4Nb34d5qbB1Phs1FrVdGeoidh6SLRE5wnnNjb+4Wuv/7uPfJpvrXN3RSHyl04ef+rgXf/g1TdWx+Nbzm+LO/P00l/jk4/6TetT2pp+6ohh2g0JzVpmO58FG2zn2AJNgbvnk7TPBsQYvIFgRU7333P46aeeeOyxR4te78KFCy+88IPXXj89Kr1XBCMlMlUEEBvi7iMEm4yEyeVBA0AU78AGM4tuXOpDZKs9eSDuZApQrWPtKohBDKa4Pkqhns5a+de3yTbXbNCAuFNl0ryTpue6qwTok/QlG0hWkGREzGBqbnVGFohATE5EOEb9DQSTFAMi+YoJkzCYwARmikZYVVWGsSKoqcUFe2ZhyStxmXFgrkg2Vd/Lsv0h/O7LLy/QUR06dOjQocPtREdAd+jQoUOHjw+ceSoLdmUZ5NrGWq84IOI4jC0ErUYA+ktLo7Jav75eZBIJTCIhsGMmxyLiREIIrqqCqsGIqCoryqW3ZxDpKCcuaKjKSk195UejoYgYYTQa91T3EPmAUnlcrj98/2FlXq/eOrs6Wh15qbfRTigOTHYHW1BflgSAidmBYEmhjBhusNJQAkiGqlNPrBN9FqVH1JirmjpxIpykVECeZUQUgxCaaVJjAWoKEBNlWUZEqhqSFjjxEVVVaggwOOEsz4hQVWwVmQZLj8TU5ijm7Lym+rJpjqK55ieIpI4OCBCIRRozkCZlTbPFx+gMdRMSEYRToxpIuFHAWZvaoMlDPrOLTiUAQghEhFpWPE2wEMVggzAYsTgzMw3RfoRlWsFdX0Ajx6YZkuHmtc/W5uwyXkgBHe6g3wG1fu4KazdTBBM9s4Ab8ouXr8wriwBbHY/evX79xMouGt6+kycO3PXdjy7N1qdeIJihxadL+bhRhvA/vfLqpdEIczja7fYc2JYXC+H85uY33n//S8eP75ryX3nggVdXVze8v6H8d8RsVT8GQpqIakvtmSWg9G1t3bvm1OXFy5f/l9de/7cf/lR2J3XQESdWVv7GU0/89z985f31m43jtp0T+fQArxdaZr6edW/s2Cu7eXbcEFr7U+Z/fAPDI25dIlNiZEx7VwYPPXD80Ucefvjhhwz01pl3v/O9F8+f/3BU+spbMITI7oagwRMzSA0etV/TlqoQkp1U+igQlMhqybqlWYBbbDJAnNJPAgU0V4a6t6gOexunm9p5I+6taZH7VHcdpV6wnGRF8h67gl0hImZsJnHBxZRikAQRojSNBo0BE4nZmXBIO6vImxE0VKUQnBORaGkN1QBTR+QcZ3nu2GWSu6zns97aeOQhpTc39IdyfCTZwh3VoUOHDh063DZ0BHSHDh06dPj48NO/8Pzv/tKXS80Iuj4aZVev7l1ZkXJo46EGL+KqcuzHVVWWWqXNti4vSMRUiTkxuQQIV1WpMJdllQUQlpYGBESPDjPLiyIyucWo5zIHw+bmBsyEEYKNSt0Yh6WVg/lgcL2q8Ma50bnVsh1ACNMvzKCmZtHkwokTYmGOPhswUw1mBmK0wnlF5TUBPgSrpbVNgKPoRwmDmWgNU20R0NPP8hZjHWncsFt5771v5LohFgEwZywszkWHbF81uubWU3r7gX0OmTOHQ5i4PSfPixYJMq1CnbgVp1hhlExCZghes4bIhhFhWsQGAixR20RgIoA06Zhtet87TfjxJvhiY0M8LR5sfDmpVdEtl3praLO3C53gFkx3k7ihzGepnEf371/JdqEq1OwHl6/skOD7ly7vSkADePbwwWkC+kcUoxD+/iuvnlm73habTq08AFta8pZG1fPvn3364MFd3Y1X8uxnHzj5K2+8eStlfeIQat+bbuar8cKlS//tePxXP/3wwd4u1jG3jpU8+48ff+zvvvTy+c3N25frdhfeXpJBbZ/c5qNb507NZbsOv4XGp5nRIqtl23Zam0BPt3aYMrB/794T9x198jOP3X/vsX6v99Z751574/QbZ96pxsEHUyNNpG/0xbAUaDctctZa6qmi5gnGrS61Xk4lcs3mJCIikjphWiimNh9dTyXRBQTJWSty0Fona7TPlq4vTZ2UsfQ5W3ZFAclADkxQmPJkNTRS5gzA1IKm6MjCZMI1Fw0J0YhbLXhhUsCBDMiYhVkYmXCeSZ5J5nLniqxYul76IFnlw8awKoRWSv/br7y0ez926NChQ4cOtxsdAd2hQ4cOHT5WfOFv/eY//s9/rjQsWXV+dfXq9bXMVDdWV/pFv+htjHyWFU7ccHNTfWAiF8wI46qMDhVOXFbk4tzVq1fVbLA8GA6HROScOBEz82UV2d6lpaWiKLIsi4+Rg6W+Bq/eEywoKo/g+sv79y8fOODDn1y+vHp5hGDx4S89Ps5CTX2ouBJmx9zrL6tqVYUQQqSYiyIHoap8NMqovM/z3DkXowtGUR8zZ3nmvY9eFlRre9XUNBKzBoBrGTJFCw8mUw1BY6VEJKRQhwDAzFElzMzQkKw/RFiVqqrFMO8YwcqSP8bk+bwBUWwOmy+nU0yxEhNChIhR66NrC+wZ85GpI3OyNjUPi84nNSHdtBUQZdiUZHB1zEZoIxo0M6NG/117eKB+U1clJW7Ic7SOL4Y54j+vC52+jVRzwaJ3SHZzCtApyfEi/hun19auV+UOCV68dOlnT57YNZ9H9+9fzrL1qont1pYST2qFen2ifeRjw8Xh8H9+5dWLw2HDbDXrHC2xZNogMDOcGpeXxYqaJFOzX3njzb/+1JO7Okv8xJEjf/LhR29cvbpYEXVJCzjNbG35OwSuV4/qxbUdxO+pYltlwO9cv/7L33vhS8fv/+fvOSq7NdotYilz//6jD//t7780CoubuS9cpa0Jae5r2i7POZtdbjYZJYXvTiNgh/HBTFrnUN9bjZmE7fj99372mSc/8+jDZVW9/c773/7O999+/3zpVY2MGEwEY0ABZgZEQzAYiWMnzAQfZr5XBAbI2nQ9JmR0TErEwk5VgwYAwiziAKiphmAAEQlLVB3Hq27006aqIWjwQYNhSvg8Mxdw+k8DKZalKFicgg1QNVNLA94MpqakMBJTMw1BvaoCJtFfIy7FMokwE5h50Cvi1efOFXnR6+W9PM8zESJhCIOYyRXrw3K98hWsguvt7Y+urf16Z/3coUOHDh0+IXQEdIcOHTp0+LhRGiSMN4abnBXDoWamYVhubo4yuhaMRPLMZUwIPlRV1RsMsjy3RD9ibCUNR0xkZkxUbowZILLh+qYIAajKCgZm1hC4Fk0TkYgQWQxmR0TOkaFcyfOH7t7/Zx57sBz5P3j53SubZSDyarOuCLW7gME0hGpcFlnRKwoAWpgPvWiWIS4306qqmMXMyrJ0zjknluwdSVVBiOEK2wS0iCQb6MikWr1lF5MnWQWZ1eeaCTPnORGpmaqKCAGqyhLj7IFcJHLMV5WGGMNwwkG39WINC7stLbLNJxPiuDHoAGo2Nwm6GjMNS/KzSYTDCc07RaPMlAECJYMSSxnOGO+SUlNqytA0Pq8nuRpugPa7KcxR3xms0oUIqb5r/zE2xbcurqKlJnzj7Fk7oBFJzgjK087xXOSJu+7aNZeXav+NOqNpzgf4aDR+f33jvuVdBLxC9LlDB7957vx0ZSZKzlZFrSGU7qB/yTQM+PbFi//XmbeH00EjW4N+UrFp9nmmqosvLUwGw/vr67/7wQc/de+9u57286ce/OXvfb9SXZx3bbXhzPCrj05she54c3NqLppt0tnSJwO1naxp53Hw/+jM279//sJP33fv5w4fcneShj7c73/5xPGvnj5zm/Kj5sfWw9PvP+b1lxtGMm6Pkt2Jw7vF6A3C2Ldn+eTxY09+5rETx49fu7755um3X/jBy2cvXtoYluxyi37G0GZJmJgcMZzE6HtplYKY4kJjzBwxkABpM9U0U2pLGE5EEpdulRC9teJScT1XEIiZo3sU0tJlDKxroapMg0X/6Gn2mSbf/KR9ZkCIcna5CBuZqVfVEALUoJkJmar6ODeKiKQQB+ocRMSxCIsQC0OYnBMmcsL9Xs8JC8O5zIk44cIhE0SNuAYYsYGvV9XYeFyV8uAjurr6W3/07TvS0x06dOjQocMC6AjoDh06dOjwceMrz33tq3/jCzDRDW+EkfdUWaUB5WYMb88kg14Rgt/c3OwvLxe9fl7kzMJE6kN0rhgM+sxSjSuXCTONqs06Lp/G50bvKyJCzVaKExFhRyAwwzGHUIro8mDw+Imj5Ti8d/Gav3j1ehkUQWeJFkJtTGoheDVfVWbKxMJMUcFKBOIYYDAqoKNgNwmYiQB4763JrhYaxwCGZqZmUu+ejrbHFmW60Qk68s4iAEIIUpsvhxCUyDlXH2cmaAhmLE6YpRIpR6PGM3qODrqmblp0xnSCeuvxxHNgyvSZZw7ShHqe6N3qz+Yxqo1CuU02NZkxmaopiGCqUJ1otCO70Xg51yGnom6SSVDL2eO/6ctrM7a3gkaiSVP1B8r50QVnsb8othzbVWe6SIJd0SJj5mX91IEDuexuY/3i5cvb1a3J+oXLl3cloAE8e/jQNAG9XcYfNy6Pxv/wjTfOrK1NDV/byj4DDSXdOnIraJYWfuvd9548cOBIv79z+sP9/s/cf99vvvPuwuzk1gFwe74a3/noo19/+51ZF90tawZxo4Rjypn7TuZ5WFu9qDNzIqYo6DmwD4fDX3nzzd98550fP3z4c4cPHdvNxuSm8eeOHvn98+cvbA5vOadF2Oc0cyyS0yeIZpmTbGpHESWNcNizvHz/vUc/+9RnTp44nufFD1974/svv/riD98AZ5LluZBatJ5K3h8GEMUNP0zExhw/BXE9OpoJlqZnqdbuF5ukUsTgCmkK03rJsJki6zAPKSJuUIWaBR+qChZgM5tcUtbUekMAgzKwxFyS21Yo1aupkakakUUrEmZiMxIWJjJxjqKLs2NxJE7ICWVORNgJF1nuhCX+AUGAqSNlkBmZAiResb6+PmYaDe265/75D/Kjx25Hx3bo0KFDhw43iY6A7tChQ4cOnwC+8rd/96t/7afXZaXwq0TIe0XPLesoZ9NqXFXleHO4GXxVlqVf183x0EnOzEwEg2N2IuPxiFmyzDETCzvHke3Nsiy6VjjnmJhqPqXy3sNDYTBhqPB4XAYbjkfjvgweOHbgc4/eH4AfvnORrN6h21JvpadmAGaKMNzc/PDDDxOznPjl5DjRbB1PqQ2xPgCqqgJRnmVJ76wqIlGmHUIIqnmeM1FzPBbLwjH3RocY6WZVLcsyirtjgL4sy0SYCEGYDEzEAx6PRutAOR6HyQP4FsqmNsesfZtpWjA84Za32mXMOwKOTdE6YluSNbEZazfQVg5o03imABmck9hoM47STd8wc+QoVUMMkGhmUIuhm2CtQpK9STvYl1HNnE+46cUUttPS44kSe6NaKBxcT6QnUu/fnyluu9Jnj7fqcKPOG7MlNu8X8d94f3398mi0JSOqs0ovXrh06UvH7981txMry0cG/YuJxWvz4wZQS+ROTQHzLuH2oxD+4Pr1elhMlhmmA6C1D7ZhaDfrDfCCkwsGUKn+6htv/rUnn9j1/C/ce+93Prp0bmPByHg283pray5o4zCDSvXqeLxjkhkNr+0w4Lfes7YcsnnpzAzXyvL5s2efP3v2QK/38L69p/buvW9p6chgcBvdOZjoJ4/d86tvnr7ZDGj65ZZ1uPSbZhPPEtZz7sbtj3btylp7fvPfqVk75rps4kgTW5pplB469cAzT37mqScfv7p69cUf/OBb3/7Ti5evuqIfjLzCb45gRtA4BRgBZoGjBjlaS9UBb5k4vamHEDGhNYsZkua4fWVEBBYn7ASAhuB9iKeKc7GtQuXjzKumFtSCh2q0qyJYqwSKR7Z0DBgmxBmJr6pxVSnSGA2EGHSQJRMihmWOMsd55pyQMMg8M5xQFmNOAE7YOc6cZI4dMwmElEEwhYFMSYlIYGTElBejcTUKXHrdJO6JDNfWf+MPvnbT3dqhQ4cOHTrcOjoCukOHDh06fDL4yt/9nf/uF//qe8uPP3T1WwqqjPrL+0V9lo1CmcO8afDBj33wqj5UpJGnNI9aW8zEJYskgpcIwpLneaRuRYSJGSROmFlNiVmEiUiNghmBhZjMHOm+5eyZR+8f+XJtfe3CtfH1So1Irf0k3t6cbqHym+sbLsvyPC96WaRAWVxkraMm2pKbRnqkN1N2QiDiSCkjhHhJ5MQRMwXvnBPh5gm5UXM7cUSkarWjCDKXsYgm1pKC+shEM5Oa+soDxkRZlmVZLpJtrK+PRsOyLKNAuLVNuIZpInIjAUEA2iRyTa7NSNniESIW1qBmlvyoWxxKYqinDkWVdx3badqaM0ZijKpwq42zCWBOgZhgoEQOpz3OQG1cAoCMWZpSkFLQRJHanDnDxt9uGnN1F/ZtgmNLS6fX1m65wBti03a52pU8+/S+fbvm8tKc8INzqnFhc3h+c/PoYLBrhj92+NDX33lvkTzb+vlds71FLGfZ54/e/c0Pzm+pzI0WfUtVPb229vvnzv/5e47unEyI/spDp/7rF168lbLuPOY2xZ1VuV8ejf7wwugPL1wE4IiODAYHe739RXFXURzoFXf1egd7vYG7yYejZw4d/D9Pv+0X2/ewLdrsc+tQ68XNDSFq1vVmNOlTidICpFmbu229muPXP4fRpsYNI96vkxmSKqBEJsJ37d9379HDTz/9xPH7772+fv3V19984QevnD13YVgGzgs1MoUGZWamJEyOpZtqCDBEXXRc/CX1lohdaoql5mIAsjg5xRjFAExBDBCgZoECIUY2jIJmJQshtlSMy0BJh63JcCO1TrNeEqehqSaLwmdH5Fh6LDk5URMguW7BmAlEQpRz5hIBzVnGWSaOSdhgYFJmY1JG3ApkZAYLaf7S5LOTZ8mKA8RmpCSutzTyYWgojSrjotcbj0bPf//7C42UDh06dOjQ4Y6hI6A7dOjQocMnhiu94/dcfzUrKy0yT2IsxWCJfeHUMxRQg15b39wYjirvawkUYtQ/EQeFBi/OERB8GUMGiTRB/4SJmDjLXJa5NhAtMkTEOZYsqC9EHn3g7tF48+rqperM6vjqaGxo9uxGQ8m2C6qaalmKiHMy6PcIrGqSZQaE4F2WgziEoDUBHTSEEMS5SJ47J0SkQUMIZpY555yFIM45EXHivPfe+1SigYWFHUCqaqpm1u8Pev0+E4cQfPCqAWRMpGohBBiZKTNJ5sQ55zIDKVAFtaCA0oR/TTDTWUaCJO4bnkJN2DY2GGpGUccdgmkgieQ7Ep/cuMc2PAVR7Vgxj80AGvcSax71mRmt3fuE6GuiaoiJQQYLqpETYE5aP7M6PFS0n9a0P7oVi7DeMT1Vx4bbvFEubCr91XJRAvq+5eVdCej2AshuqXbFDlLThM8dOrRryDsAy1n2k8eOzeS1taoEbC6mB3/20KF/8s57zVhpfTIZndO69EX5uDi0FrmoufjJY8d+/9wFnZKQzlzobDPM7bJbI8vpH7/z7uN37T/Q6+2c7uTKyp+/555bKuq2YhteeS7TejME9Nb85x5p5+7Nzm1snNvYmE5GB3r9EyvLp/buefLAXXvzfPE69EQ+vW/vy1dWb6zqs9iRfZ5DGi+YZ2v3R8zJIqM7fxmgWROcugXSVnHz1AFKsuRI+sYJW0HGIBBUNcaHHQz6J07c+/kf/+wDJ09o0BdeeOlPv//iq6+dVgAsKMeAwAAFACNoiD7LRCwGM4ToyGKmDCGChhDj9SUvDm2YaDALiCxUhqiUFoJpCMSIidUboDAGM4mL2Ybk804kAouRcK2ZfYjAaWKJonszM66buFl/cEwFSyF5wZITi8IRZcIczxQigIkLFgExTAROOGMWBpNx8hVRi3EOAQNpMCUEYpAliTeTcF5kObOUlVYKJfHB1sZVZVSaxwOnaHX169/61uLDpUOHDh06dLhD6AjoDh06dOjwieG555776n/4FyzP2GUsrMxFvz+QpVxLgg++LKtxXvT2VH5jGC2eyfuQyFk1731ZIs8yEIL6yIiOx6OoBRbJjMXIqmGJobmoPkbt0QGwOBIBsRQFFz3x1X2H9v6Ln39Gszfo9IV3L15TMwIxsRm0Ft0C2lC3VVVubhKAzGXEHMajEBXKLCAOmnyXJVo8R2UcEQAXtcrM5XhclpXLHNfsKrNkznnvfZiOdQYmYjMFICIbG5vRDzqaeZRVCZjLXHy2jXbYZmowVdNgBCIWl+ehqtSb3VhQPmsxsxPhacPgqpkH1HuZyjoLAAAgAElEQVRT9fVO71jpLUalBOIZAqUx3Ey6MlMLGkKo4z6BmY3Y+2giYkRIQQmjiq25Xk0cuqaLMw0Bpmh0cKYNdZlCNDY7otFc2W0TYH40HC2Y8sG9e7557twOCXbThd6KNHI+Pndod/8NALuqcW8UB3rFg3v3vHXtGhLR3NCGiXpGUsA3VNyiI/ncxsZ/+b0XCuGBywoRIVLTUi1j/sWnn3S8i3XJ/qL48SOH//DCxW1oZbPpXpqu/OTwrQ0vK4P/tbfe+o8ef3zXpF86cfy11VskQ28Pthm9N0mmzsXW/G/uCGCXR8PLo+F3P7r01bfOPLJ/3xfvv+/knpUFq/HAnpUbI6An8v36VRMmrxbzYvor0DLonhld8+n7bcZbunnXe1CwtSNsKrbeLSE68DMTswwG/Wc/98xnPvPIpx964P333nv9jTe/+72XP7p8GUJEbNFQIgqIRRSEuBHJEoU9NaHEHTEU52QCEZMQEWoyOAS1uFYZYwkawJQ8o+N/gCWaSpPVLDm0UYtTvV5FGlQtwDTagZgpNcub0+uUsXABeuIGWZGLZMTOiFnFIFDidMuKfhkc3Z+hrMwKVqKouSYlaLrjxdoxx3iE7JilnuMMQanyBthw7EtFxajGwTse+nJ1rIML57O7b/NdukOHDh06dLg5dAR0hw4dOnT4JPGV/+GbX/2FLzojJZATwPorK3k1ND9SQeYIkvXV8iKPj6Fq5quoDkbwoazKGH+n3yuC9+pDlQygM4BUrfKVaTBTXyXT4SzLJUYGFEfEakZZLnkueU7F4PCewUP3HVrbGK1eXbteYRwAmDVPtADAhLhT10II5XgMszwvXJaFOuBh2rgLeFUz05opjoG0zGBmgZmAyvugASFuUY6ErYYQQghqJtHKA6YhxkqSyEq7zPkQmCiaWppZWY5BlBdZLFpEiMzMggY1wEiEQZAsS5yC93ET88Id1XAeszxFfELWRP4mMXGbJZh1FDWdtsluye1Q65Oj1UeSTmt0DKmLiDS4mikxojKdo4G1NdRMnW6idG5dhlmKG2nTJs+3KyphjXMbGyEJ3XbBI/v2MZHO7445e+HnJbid7PPhfv/EyqKk223Hjx8+FAnoubDp6906IHeAAaOgozDGNCv6px999BNHjux6+hfuPfZHFy5iwixvxW4rBbcDr65e/aOLF3etcE/kqYMH73RldsWO3TOXg/442nBHWLoNgV5ZvfrK6tWfuvfYl08eX2Sc3UyQw60c9LbHrb7dNscb7CAxp6mFw/poO5NtBvQN94JRI3yePt8gQs65Q4fuuu/+ez/zmceOHDm0tr7x2punf/DK6+c+vBQ0uF6hILU4ezJIiB3UYCBLG3HM0l6WWunMJELEHEPyphIpWkIBgPfRqqt23jBihqmGQFEZbSYiIhzF3WamIcTNQJO7jJkamRkFqgXPStH0yTAz5VCqOjmgYNcTcSAxE1NWE7Iodo7WW0TERgIwwGYCExgDYqmbKfLrcfGZmVjAzliMREFmaiGYqoaKEcxIwZT3vGpFviyhm+Ugk81ra8//f39wo13ZoUOHDh063Al0BHSHDh06dPiE8ZW/81u/8Z/+xd6610K9BphJlnk/csz93qAyywy9XlGWpQ/eORd88N7neQGQ974sx2aa5dlwc3NzY9PMmEXYjcfj4ebmaDgSESbyvvQh7tRVJ8JEYmrG3ofy+oY3c0WGfGD50r0H9ly/9+D5c+d0zZdBgxnAgAAwKKAAJx20WfA29EHVCkBcJs4RUTAYiGI8QTNOrhTWjuWnqqX3LFxkPSIyNQ0hcw5A5b0RhCXLXDwlqAIkLChLVWWOj9xQDWYGghExE4sEROF1QHqgNmZhlsp7AFnmiEDECtMABL0hloGIhHmGMKp3R5OJUHr6p2iCEdEQ3Qvw3TZhr22GHl6wihMhc2IrSNJrWKye1dcyzX5ZzUDXKltggQrYjCixDW92YXNzEU6q79yj+/e/fGWrnzIaTr+u5PwEtxW0SPjBO4enDx742ukzlWqLeGvsLKYu9kapyinhdOv4//vBuUUI6CP9/jOHDnz3o0tbP2pVjFpk4Zw63yhoMrom1f+/z7z96P79N2QQsVMJdwxN5VsNPiPU3cpBz1fyUvoiWOvjOSnndfHsMJmXFWhKnD7FBT9/9gPH/BeP37fTpQIADvSKXdNM15mmr6A10tGsyAELy/y3K2YKc/TOFjeDTCejmxgbEw56ukAhWuoXjzz8qT/zEz9299HDly5f/vYLL37/hR+cu3Ax7/UcsxH5GOfPACMiERYLGmMAIHk0a5xXo0FTDDkQCeY4y4/GYzUTEeccAex9k6AJHGFmIQRmBlGICZq9RKoWfPKAikugZsEHX6ml9UxADWZG00ubE3coEuKcOGcumJ2RBGUNsEAAM2UZM4HjRiAjELsYbIEgBCa4pKGOOTIZI4YxzDJiAUmAwISVg/e+ClUZLJTqVYMt791bCJTZEzaGZb6ynF1ff/6VV260Ezt06NChQ4c7hI6A7tChQ4cOnzyyUnW5b8iGvrqytnpwZV/RX9bx+sbGpmSZyzJxzjGpZqoKESpyl+VmKMuSTIP3bBj0+v28iPpiU1seDKrl5T3DFWKY6uZoqDAiBhCCr8rSggKW5y4rcjV41aAh+FEudHA5//TJo+Hty2W5PjLyBm1REg3nGB+MVS0E773vDQZ5XjCLD0EBFokPqcSspho0xuurIzJZlgUATCzCzY5rVXMhcAqyWD9mhwAQs4hz8eriM3WK1GeWZ46FnZMQIwESIQU+NAIxS57niQF3mWa+ZFRlGeChN6CDNrOgOqU5Jap9Myb0OswmgbjqvLmxONiq6G1xwAYwk6mpapu4JyInEgNJgUDR+jPq47j2o7bkN821zanGSFWGuvBE5TV8dGR4CNFrulFk3wDvPZ1wlv569/r1BUWR/9zdd29DQM/kf+cwaYEF/TfuEPrOfebAXd/96FKbxZ1L4960UHbmxHMbG69dvbpI0MV/6d57v/vR5W2ybKraHLoN/TX3Gje9/+rp0//eI4/cev47tuJ2jP3iWTf60CaHm+y0GanplqxS/jbns9kS52W1dY1n6vb02++f/bNHj+zK+C9n2c4JpkHt39Nafmp9TlsPbZNyOsHWzSoAFu+A9jrctmgmrtmMidksRF+MXpEfOXTw6aef+NSnTu3ft//M6XffOnPmldff3BxWebFEIj4EryHaYkhNfKspMRiJIAYADwJS0GEzNRVmTiF/NZhlmcTKxPCBHMMQkwUNMUSERuGypd0mxFALvvIppmGMOkBwFM2mVYN6X3lfmsYIhCFOU7OTZs0+MygzKkh6JDlJBiMYEZg4Y3ZCwnGfkxEsLnpQvBwQYtRkl9TcBKMmUAFZ6YNZUEOou5JiUERVJ85lGQpXDAYBVoKD1+KRR/xHH/36H//Jgr3doUOHDh06fAzoCOgOHTp06PDJ44t/7xtff+7nmZVI1yuS9WtH9u6hrO83NwVgokzYxVB+HswsTgBWVXKO8twnSw1mYrX4z5hEg/b7fZgG9VmRxzQhhLIsx6NRqDxALsuNOKhtDkcgIyi03NejB+85uDlU73H+2uYwmIcqiAgEotbG2+j9oKree1UjYuccMRtRJKABkETVlaoGEEnNGhsyMyND5lLgRI0qr6BUa7YiixxCiApoZmkEXEQU3TmChuhjSRwl1zEKn0UGFqglY0BQjedkwmNxJY/LsjQNyVNkFpOwS6h/mZlNwixF5nfLRvEJGVGfyROWZMKzUGrGqUBYBCIGKyXambSO/sTMUA2UhMzM0RG7Jr5rHXZyTaX4gG+NiDA2ZpKWTVtzNGrDG4TN029O4dXVq5+/++5F8nr8rv1HBv2Lm8Ppw1uVoXccJ1dWDvf7H09Z2+HZw4ei0DgJ4mf6KrGNW5cyFsHMiSn33/vg/CIE9H3Ly4/u3//K6tXtM9+hxF1GyzRo3ttJW7xw6fL3Prr0zKFP3mTjY8csG+6YT6ys7GDbsmNWmM9ap7epF9TsB5dX/+zRXWTy+W5O4luKnss+tz9vfjXpp9b/5qWub8hR5z2VYxQ/b+FPZ9thVh+9LfHdfNSuX4yVQBaNI7JM7j5y6NSpk48/+cjK0sratbU3Xn/z9bfOnD1/kUWInCqCN68mrl5ITNtTFIh8bbpDN8udkX9FXOtURZw6zUSEANMYntYYgDCYQ/AEgigpmZkGVU6KaNW4MUpN0/2cQcRR/qzBBx+qEAKZWiR8MSsVr7+ZJECGxD73OctADmlGY4IICzMIBm17QzGREdfdyWSUPLDj3Bip/WDmvYagagomgjAVGTtHTNLLc8l7yhkEpVkwH8B04YJbbOrp0KFDhw4dPjZ0BHSHDh06dPiRwJee+7Wv/xc/d6XEAYero3HPbexbWuotrTACAQwEU2hgMmEI0Wg4VDWXuUG/IOoDUI3uycYucy4ry9LDepSpqirXYf84hBB6PVtaiiECFTQuq83xmGJon0w2x+WAcHRPnx66tz9YXn/htIaSoBVAJJm4EEJQNLuAAZip99X6+noIOhgMXJ7FCIFBFWa5c8Tk2MrSjODEResMZo5bjDNxBqiGjAUsJhbNnbMsj+Jo7z0Ruyy3JFgmJ8zMBlTe+6oSESJS06h9nqgwiaK2KyXQoGqmSoP+eDze3Ni8dn2tGo8Nk+h8LTbGQDrZr524i/bjt5lRQ4IQ0axDQsNKKIKFNlPR4vDbJwBEimRsXUfIQtSqq5PIHUTHEWNJRLKP0RoTJW0aiKWuXosOb9Rk9QdTVwpM9NFb1ZC7wLYwOOnFK6urC9pAM9FfOnHi77/y6kxzLFiDG4FiR0XrJ+u/EfHo/v3LWbZeVahXFmoNbc2g3Tw1nwZ0re1Mff/DK1cubg6PDHZn3n/qvnvbBHQ7K0y1alMQTR9ZaFTR1KCautim77525vTD+/YtZbfhj/mZ4VtjO2b25vKeKqT1ZisvT3W72ryBOnugL/JvfuqhX/re98fTgVu3q8f0gXa2zeiac/zSaPeYogs306yaedIENN3XM7eOaca5/rS+CU8XT0A9GczSzUQ067nRjN+FnDcmFUuLrCliHzEzgUxV1QOW59m+fXsef+KRxx/79L59K++/+8EPf/DaW2+9+9GVq2UZwBoHugHC7EhCUO8rEo6xAU0jNTxppjThJtWzld5bsLjAaWYVUFs+EQCEwHnGzmlQIvLRDFoteB9Xo51z8RrStilNBRh7hFi4T34bqpjEsJ20J9X/HSgDZeABZwPOChKGEQwiKZghcwwpaMaRMI+5aYoYbBxMNIgBFkyVUqBghRmbCtRUmUiyrJ/ny4Pirj2DImchy4s+F/21cbm6OQ6KamhOS7++/rWvfW23fuzQoUOHDh0+VnQEdIcOHTp0+FHBMGApcz6XrBpf2dwMAcuD3sb6VYTRUi+PEfmqqsqyrFewyxwROec0NA+cBlg0rlD1RGgeL6NoNz6mVlWlqgT4yodgBsrzoj8Y9AeDAAOoX/hhqRuluaIPluvrG6fPXTl/ZZ0Qd/36+Ow45XRpULVqPLIQfDnmrGDnqJbauuEovvY+xCdtqqnZ+Kocj2sbifRYH3wwmC8rFqYYbNCIaFinoKSYrtEYXEbr5zYBTSAQhAUEjQJpM5CGEMhJv99nkaos1QfTsIV7mSaIaCvBMmFOZoMNTs5PJ8/Qu1GYnfpntthEEyfHEuYWPTRFfDSl17RJ3AZN9Z7o2lPV2h4bkcObMOGRh0xa6RnJ4A1w0HMwCuGta9ceXkBaC+CJAweePHDgxctzHR5uCwzAvqIoQ9j0fu6nTPSjIKoVos8dOvjPzp1PzVoPw9SXM+scC2fb5lNbWcWBa7937ty/durBXTN5aO+eB/asnFm73q5aTTS3h4Ft/cJsoc53qCrNqW89JOObtbL6R2fO/FsPf2qRDHfADQzzm8EcFntLiXM1tsBigUEz5gO93r988uSvvfXWdmkWIbKbfpxbveGcr8wsRjsy4DMZbj2S1slqWpnq29PkGtB8gvrT9ura3Dbcck9uvlTTd9B6xWSR8dnKJC4mpumQNBizmCmg+/fvO3bs6KlTJx944L6il73+2utvvvn26TffXbs+LMsqVCVEwBznOACh8tFVybxXJaQlxtZ1pW9qij9bR+GzZLQxuRoy1fhV06AGH9XNhGgMAlVlJg2otGouJ3pzpK1C3kwDVFUDpelezaxmy6dajgEB5SQFS4+z/oR9TikUpmZQI8DUEpGtyWFDY1QFNWZywqrCjOgTzUzMjmGOkLEx4ITzojfoZSv9bP+eQS9jYphklhero5EJvNnS2lpZFF97+YcL9GOHDh06dOjwsaIjoDt06NChw48KvvLc137n7/wbWRjlMh75pUvXN33wVal+c70cSa/IhXk0GhVFEYMOEYuaVr5SVREXqdhoi6zqiURS9CGkHa41nWGqRMSgwErE7DIwL/lQBu+9N2BY+nyzXJKi6PeESZjLUXV9XI2CVkFrCslm4laFqgxVOR4OKSs4y0Si8pWIxkghjtQMBBInsZ4iIszxedixBFUYmDkEr2pSP5yrWvwfvUYS4WoWNCQCzIw46rkM0AlvQYhaMkrpFVEiXWtJ86IgYQM8KvUxNOE05zMr69yBnpgldHZ2Uq75ZzT8wvzkFI27Kcr55gj0kmUmxc3M9fuJDC62Rc3ZUM31tAxGDMm9YyuLuBMWSvrtix8uSEAD+Ncfeuj99fUr4/GC6W8UOdN/8Ogj/+trr7cJ6LYy9NH9+1duzMf2TuHZw4f/2bnz8XVbLXvT7PMWtEkkA/DHFy9++cTxgdv9b+P/n703DZIkyc7D3uEekZl19PRR3TNd3TM99707e2CxEEER2IUAkBQoEhBMgn5IMplImkmiTH8ImiCYbGQmQUb+kMxEkSJoRkgmkQRWEEGKWICACGAXx2K54C7mvvvu6buruuvMjAh/7+mHR0RGHlWV1dMzOwOLz2aqs+Jwf+HuGVHx+eff+5GTJ/63N2qt+vQpi8nBMaP2eRI1V97k4eKeP7px83NLR547dOjuSt5nDPv7esxa5PDz5AF714UAnhgAvv+B+69sb9VjZrKmHXXe44cN6x66+4DN4u88C0k9xDgLbaNdXQ/1OpDqmMZcX2OGEIZS6NELGaljuNKl+eyq74/7ih6Gk51WqpMx5tMjTJLOiRMPPP30E889/yyi3Lxx/eWXXz1//v2VlTXnuwqmKoBxGrLM9ychACASmqgKGNU+FTRSr1nlg2GgOrwoRKiSDZZPMXbxQg0A4tIfrtoSERCkmjCo6HRjQgBQFVMFFah55wb7DI1RiwAE6JAS5pSTDnkfH6hxshct2mBplD5bzGGoaEZqaECAgkYAYApMYIygLnGe2RGwI8fsCD1D4sATJc51Op1uyr2UF7su8QyEBae3twd9LQKYZMxkyYf2BGnRokWLFi0+CFoCukWLFi1afIzwI3/9//qDv/kXcnGAg0z89dUNT+KMb69vMmpMT5cm6SDLRUVVzcy7JE3Thbn5uIw2z3PvfbfbVVFTNVMwUAGNmigDMSNCRqaU0ACRVEHMPJEpIXOSpt0edLq5cHoY/PFjx+a7vbnUv/T2+zc3+goglc1wxc4OlWkAEEVhhJSmCRFhTIRkqipFCGZAyBzXF5sRMSJKnqmZmAVVAHCAYiYqQTUy5OWrPUAoJOqCnXPMhMxgpmrRn0SDESENCQpEAFVBFQNTNVElImQcqrOZkTBNUwIsAEIAiBw0jBFrWF1ZSdoOlciwT+KigoqN1lFTK1Arow0MQ1OlOjy2lMbVhAOAqSECEpYOGxNApEr1bMPqmirtHcnDnYANLmJIpWEj1pdu3frJRx+ZhdYEgDnv/vPnnv2fX31tsyh25ebuBgnzf/r0kyfn5xvBAwwv1eC7nX6wiVML80d73RvRFBvLH2YjrbGvdJHQ7CQcKwoRoFD7g6vXfvjkiT3LefbQweW53uWtbaimNhpfmHp6aLTq8RpnjLc5FsubQOlmXuGXTp/92c8d6NSJ2vYNtCmjF3a4nEnp7u4XgM3RBdVtszmjBbv1I9bhNEKs6cZYrrnKefknH310PS9eunWrWULjy1h3fv3L9C5rDJLhCY/dt7jn9d7s723TMYLmJEj5Ozb+rVfZaEU54+j3dRRxrhUnNs6qa/6gICQEkJAdPnL40Uce/sxnn19efiBx+Nrrb7/++pvnz1/a3OwHMwmFAYAjQDCLq31KfhapuYSlDrsRPwIylvdtAsIydwLEmUqsVhcRAyI7rpIoaHz+oWNAMFVkJiL2pY9WdKYCFSvtOOJDvvyv1j7XrU/DS0aH7IkT5x2ymeVSiAEhikoIYmSAFvXZiECGDEYATMgGDJAQOgQCdI68I+/ZO/IemdE78o4co3PgHTgmz5gm0PHQ8caQg7Kh72f5na1NAcpD8exLr964//6/e+3aR9DdLVq0aNGixX7REtAtWrRo0eLjhe//G//8t37uL4WMKIRtC6HQnmNAV4QMLSTO5UURRAjRzELQwkmRF0WWIyKgIVKapgCgQWoPB0RUMEAwJHaMBqW+GAkNo76JmJGQAhIAMR2Y7xVGhVEv9c+cOpZ6h0Bvnr927uaaAsjI6/84XWsqKoUU7Lodn3iDUqflHBsgIVc2GiXHQI4jKVp6WQIQMxJBregCVDMVQwCMF8UERGBWUuzlUWgI2pAVG0K0ba4yLSmjY6uyIJrlplEgTkzOOwModdC2q9hxinYPJhSETTXeFGnecB822Becsh0BgUDFGmRz5b4NRkRRfWcxPxNhzEgVOeyy5AabUHHZVoqgRzRtdw3bibYuVL957fqXTyzPWND9vd5/+fxzf/eNN+9k2T6j2o1jOtzp/NVnnlyem2tsa/aiAUDC7tOHP3Qt7ez4wtGjX71wYdgG90p6Ow2x7N+9cvXLJ5b39OxGgB85eeIX3n53p6D2RYt/QNzOsn967vxPzWAeMiMmJ2TuWZEjk0jD4bcXNT/CWY9+MABIaHjL+0+eevIrp90f7ErATVzV3qz68V5vlhyVN/r9PY+ZXulkCDUHPQSOHDamWR5p12bb2uhCk5rJbSjyp1/9FIZ7yq9YGrSjARF45w4ePPz4o4889+wzS0cPDrL+mbPvv/X2O+cvXtruZ0ic+sSADBGiFYUZYJkmF6x0q0B0BIRMWC1vadSJQBSzAsS5XERSleqCh3MJSBSXQKlpXhQqCh6YyABEA2G5Pio+BxC1fHpKMBWIT8AmBw3jYxQBCJGJHbInR4ZgogqqWpgxUqS0ARA5GmQBIzpEBnAADtAZuEhAgzGi9+wdJ955T84hM0VKmgmIgZ05Ns+WcGA0MAoBjFiNVtY3+mI5hm6R3nz0oaNnLkztzhYtWrRo0eK7jpaAbtGiRYsWHzv80M/809/4mR/PTI1csLwv0ku6hKQhd4lXKbJs0Ov2mJxpCIVk/WxNbiOi8y5NO3meDwYDFSVEZnbsmBkYiZkYnHMiWhQZoovuFhDlSC6JmfqyPCdwvW6HssJCLpKdXDpw9Mjh1DMQXru9iaK5WQBTqN9KrWFWiiBBTPsqSeodd4KEyJ8wMwIBkpoaAMYPZt57UxMRhw4A1Myxi74Z8X2aiCRIngc3XGSMACAiqiBg3jkqZYA2bjxrAGBRglXqxAANLJZQhABmTESEzjtECoghgImM8w8jskUcqWBEPQk1ZYA1iYxgE6TeeH6tUUqkCWICQFNDKs2vTVWDxkKQsEweFamE8kOtGaxCj7q25oWMf5jguPbg32z0iCEHPXbev3z//T/9wP3JzBrV5bm5n37h0//nO+++fefOB+egPdGXl4//WyeXp4lkRwp/4fDh2YP8CPA9S0u/duGC4egQa5B1ZrAvX4thB1cnjol/7+TZH9+8NUsaxs8cObzU7dzsDyZUrKOM4UiN47tniXdMLDwRPADYN65e/fzSkccPHNhH2RMVTYuuGs/WbKV9NfjuB09OXO0ErFwXxs4FAKgV0ABAiD/1+GP393r/7Pz5oDptLmCHKYOJa6wMgcEj/4dPPjFLlOc2Nmc4qhnJThx0za4PaVUAaOR1re+09QU0zq208vW1QXnPbiYPxD0afrLlRilvRIhSYCLDkoDG3lz36aeeev75Z5968vFr1y+/d+b0t//1t2/cWt3ezjrpXORWtTTet0KCqCKiY8/MppYXRVEEcszEzMzkaEoaRlRVAENE9g6JYqJds0pHHYtHRABmNgQ11crQykxREKvvULymyEYbYyGFagAtrTnQ6gLrXqkDQULyxJEutiCiBgZiAmAKpSMIoWNiF4XMDA6RwRgwQXIAzsCjeTBH6pzznlPvnEfnKHp/ESORISmQIVppLqUSjAQZUDc31jeDBsMsJT8XAI68CC0B3aJFixYtPqZoCegWLVq0aPFxxI/+3K/8k5/5cQdZRg4UAlBn7gCEQccTSBD2JiYmZKSqoIBGaZL4xEuQfrG9DRaTEyJgkiTsWFSicJi9S3yS+mQry0wBAZ1PvE8UgpqigXceAIt+jmApoQMM+bYzfvLkUj8rslC8fvba1dtbJftc6nEnqRYxsX5/wyCkaSdJPGG0tEQAJObI0kZqgIhUQlEUaZIgkoRAzESoamYaDzBmzw4wWnqQqqqoeZeqGVjiPBJFYhbAuPS+1BAkSp+TXg+RREsGVk0ilR0Z8JIfJ/I+ybNssN3f3FiX0EioNZGccIQXmyAyEEe5ioldo1uGjPbEvlg6AgAzlYvJkYwQuT4EENGQIt9laoxkgBbXrcdjrMG9VHR0/GWUuRmvfVcCrckoxuudrhvfKIqvX736wyf29naocSBJ/ovnn/tX169/9cLFO7Maeo7TeQnR548u/bkHTxxM01nO//zRmdIP/vKZs6+t3q4Js8YFD7fAGFkzGt+//dCDs5C8hzvpo4uLp9fWayuHSRJ0xpx+dRiNErD5oT7kdy5fmcuH0okAACAASURBVCU2QvyhE8u/+N6ZRuHjrhswTE44EvyMoY7GO+Wqa4sIA/tH7733M5/9bEI0paw9sMsQt0bXNWu8a0x+O3DmJtmxqITHr/oHl48/e+jgV86cefv2nYkTRmJodJBVWxpqa8Oec3/56adOjCwdmA41e+fO2l1dyy4Y+xqNtF51E8PGwc3Js3i5ZQvbbl1nYLrz3lHxtAhEQa+VGQs0BOdoYX5uefn4w6cefurppzvdzjtnzrz11hvnzp+9uXrHgLq9OURniHHNipmJGBoxoJqFIoQ8iCgAEJKJipqKKsnY8yJKjLG026Asy9QgTkxizNYbH5cRosgEgEWRGyKRxCas18eUuQrBUONqIlEpovVz1cLNphxtsrhJzVQUlFQBAI0ScoxYmmwQEiEzMROTkSmqMoEjdAQO0CEkTI7AIXnvvXM+Kb21mCjOyKrGNMomBmqKZOgJnTdO72z019VydkXQxbWt9aMLv/B739mtH1u0aNGiRYvvKloCukWLFi1afEzxEz/3K1/92R9ZclsrxWLfMEFauO+Q18BSYJrmg0zFmFyWZYho5rx3jkmCqEh8K4yv3KoanSGhkpQ57ztpJ1KvYJimqffF0E4YGRE1BOfZRVdLzcHoyPzc0w8fA47Zg65dXdsysHrpb0RFR8eapMj6BooIHSJOHAKqgRo4ZiSKK5ARkR0rEQA69mXSxEgkoRgwAMRfCY0ovmiTiChpXEFsZs5x1IVFMpiJyiXCQISkqo5dlasvaqiopoKtfBNXInLeESIBqshgMCiyWZyIqyZoNkXdBji+a1ceZBwYVz43DGjBDDDyFENBaDwgUvDVcVAamoxKSOPa9NjscaeNHTMRwl6Sz/qA5s9x/ObFS184evS+JNm1qPFyv+/Ysc8vLX3n5q1vXr92Zm19hoYzAPDETx+873NLRz516ODsiuaFxD89g8mAmv3rGze3QlHFOEZAA5Suu+PXAo2R9O2bN2cheQHgC0ePnl5bn+XIe4VLm5un19YfO7C34e8Xjy79+oVLa/mOtr93R6zeHW72B1+9cOHHH3747k7feZQ3xdH3/IJmYp9T5kx2S+7np9HuR7vdv/bcc2/fvvO1K1feWF2denWj8uMpeOHI4Z945OFDs83fvHNnbX9JCHeOZoeN8eZV8sl3U9oekw17FVXe1G2Y58/UVBPPBxYXlpcfeOyxx049/HBvbu76zRtvvf3O2XNnV1duhaDOeyYWNRMBEWYyAxGrbgvRScpElIjYsZqYGqAG1bgbo0JZTURVlB0jERiIipkhM3MkoBUAmEjBTFVF41NOVQFAG+MkEtAQKzJDs0hAg0X2eYp2v759xdSJDtAheSAHSAYOiREckCd2RATGZR5kY0KuxjrG7YgOgQkcAjljRkfsYsJBRgBQA6qmdg0w/hc11UBk5MB3N7azbYQCXZHD8T98c+Pk0t95+dzO/duiRYsWLVp899ES0C1atGjR4uOLOZdtaTf1FpRygiRNCNJE8pQxpANQIPJbW1tFniGhaBAJRMicIJFK5D8py/um2ul0ASBIyPN8e7C5cWctSTpMzhTyQU5ERVG4xKedDiI557x3ziEagYpHZLIsbJ84fOD+4ycUENDWXjsnhYXGi2qTTYmUqQYpbLBlqmaIlCYpARR5EQNTNbPIKXNMmCQSFcmmaACgpohIRKVhBiKzI0QRoehwyawqIYiIqUoIoaZ344lExOyYIc+yIgQRSVPvvSdiNRMtFWdMrFIURcizPHE+SToHDnpaW1/L71RasBEx5jhGsoKVyQOhKY2exm/NwkRPyqUBAEwRkaNNdlR9ixiAcy4mV5QQDIDIVXxzlECbRb+V0XrLZfblovBRgeEu0Y/uqiwRdsRA5Cunz/zVZ57e85LH4Im+eOzoF48d3SyK02trFze3bg76twfZQKRQTZg7zF3HHXaH0vTE/Nzy3Nyxbnd83foM+NyRpVnOendtrWKfYcLFop6AmZTNDiloA3j79u1+CN0ZEjN+5sjhr5w5Kyq15ndajbOinmywnTLRgRng165cmYWAdkRfXj7+K+fOwo5C2hHifdQ3Y9ZQYcpV10boIzV+7f3Lnz1y5NTCwizlN7DHhEEzqH3Jn08tLPzko4/sXvUu+xzRvHMPzPXevbP2S6dPT+wfxjKVgI546uB9Tx2872Z/8Nrqyhurd06vrYVK3Dqty+IvuNRNnz90+N+4/9gDvd6u8Y/gD65dn/3gceDIP8NfhwFODNiR0+uWLE8Zeh/ZvlxqdkXUCzsXHz5qYggqxcLBAydPnnzhU8+dfPDB3vz8W++898rrb7z22hsGxsRJ0lPVLJcgoqqmJZsM5UMKscwciBgfRfGubgbRYyqISkHOE7MEUVEwI0QTE5E4zWoiZhoZagBQkSreStatBmAQt480oVZO1PGDjqjIYYx8L9vXIybICbIjYnQOgM0ckUNkQEfAiGjAcfoXgADYDNSoTEAcxdHkyjwOAkDkmBwggaiKKYEBsGNmYkBEYvbsHXpmR4w+3c5lPVgOBFIc/8N3+ocXFy7dvEfd3KJFixYtWnxYaAnoFi1atGjx8cUPvvj1X33xx8C4Sx7Bbq73D/Y6Pu1lg/X5XpcAi0Lm53tBUglFVDSZxoT2GgoBNWJOvDNVIgoiZOo58ewRiYlFtF8MCBGYJYQoxIpLsBU0SRJmjonqkIg7c1oU2cb6EyeOBHkyC/rOpZtXb28KghjoGLFUmXWamuRhYNuSC7NDcoCEOQKgqAEAIXmXmVpRhKhoVlFEBAQVJaboTB1Fyt45JJQgBlELxaoqlaZMVUr/5QbdR0RMXBRFEDEzEWXOkSgWCACESEShCKZqCAUHx46JnE/mFw9kg0EIuZUKxN25s3Ez6CnGJMPmGTpZ7w6ksWPMFCFaPYsamKnE5lZVLIOYKLnixOvshfHz8Ge18n6EY7ORf3aMsHLdHiXyxs96dWXlj27c+MLRo7uXthPmvX/hyJEXjszkknEXmFGS/OrK6jTh88iWhtdBk+aruTEIBq+t3v7CDDV2nfv04UPfuXmrJgerPWMxzIQ6GBzxksDmXgR45dbKrcHgSKezZ4Hf/8Cx37x0aTuEiTBwMrB9uYXs0KqTwUN9mAL84/dO//RnXnD7nH6YtKeemHrZgZHeFQ/0evsicHfC6yurux+wCwEdsdTtfGl5+UvLy8HsZr9/bbt/a9DfDpKLZCKI4JB6zi0myZFO58T83IH9rFSIuNEfvLpXnPvERymgH613rObau4isXtoipobW63UPHzj6xBNPPPrII8vLy+ubm2+/c/qtd999//LVIs8R0EgtiJqZqplWM5MYF90gopbpB+MEIRg7ZVUVMwNAU43ksoZgqqYKgEhUUsxYztMCGmh554+RAlJ8xkSBcyOdYD0LBuWRZpGDLr04mjf9RjtU+mVwAClQl1xCzhMTAaqRmiNgBDJziBSVygAIQ5U3QnRvtpgPAUEViQwNUA3LQMwAzBExk3fsHDORaUDSWKCZFQootJblAVAKvXH8HXthYenl9Rfv+UBo0aJFixYt7jVaArpFixYtWnys8WMv/upvvPiTQKpkorKZZ445dalLEkeIHFTVBwkFMRMxi4iEEETMm1WssKkVRQGG6DEpmU8ysxBCCMLEhFGGDGCipkGKQZ5nmSNmQAA0Ik5ECt3oBzi0dOLJk0vrm5t5XvT7g80gmZg2yRlsiAoNNEguWZ4VpbQ67SCiGUQCGhGlKCRoCIJREBU9LgFMLcqcEUFEJQR2DgktaqejXaaZqXIl/kWkSh1ZImZiDKKRjM7zAsCQ4htvyRMiogUFM2TSoELinGPmTreHyEVOoRhEdfZe3RXf8JsURi0vhuYLfQxsz96Pa45Ha0ADhIrMMDAzJeSYinCnhdMltVyzz9PzEJqNcBON8+8RfvG908fn5mbxk/2IcbTbnUU5awCv3lqZpUAsJeXVaRN45dbKLAQ0AHzP0aXv3Lw1y5EfBGMy4K9fufrvPvLwnmelzD9w/IFfu3hprLB7HNxeqOu7srX9mxcv/fmHHrzbYnYf7fsl/O8N8uiuO6Xucng5nNX52iHeK1p8DP/s3Hn9gP7Y4yi/QHuXOn6HjI1lpeZ+1qDKr2zzhlt+bBj0x1yyZgaEc3O9Y0tHHn3w5BOPP37s2DE1vHTp8iuvvXb5ytXt/oCQy9wIWnO5cXqUkBjAVHU4W4pRi2yGqkjxAVfqtxGZXOSnCRHJkfMaCjADrl5jSwkzlGtiTIGodO0QNdWyQeqcwaBQ0cEGDW662ZyjwnGMQmaABChF7pBLiD0xogEKgDlQKv22kSBS0IYVJR6fLBXRHtMuYCTTEZEYo481MhECEzlmF/XPGGNVEAF0xj436ve3c2RRvKHr6eqxG49f/zsvz9jLLVq0aNGixXcTLQHdokWLFi0+7vjRF3/5N/6HHwdgTjBX2RxkB5YOFRpAw/zCwsbGmmhI0iRNEnYuGwzUOQBIXAoGWZYVRVEUhZo674gIifKi6Pf7ZsbOHTp0SERExCcJO2JHqpIXGTmyuHBWg/eemTbWbgcxQ3c7qLre06eO3dlY3x5snbmyXgQZIQFqJjPqoKPGCo3ZO3aemB0DYgh1piNzjpgpUhgp+TI5IVNNshAhkiECEbL3cTkzxhXWRI4REFQBMJppChgQoXdO1fI8j07T3rsQihDU1Epzj/LlXWNOp6iGRiIRUTNmnpvrai/NBv3+1lY+eza88XxsUzwq1CakdhNAANAxdsnMDDQ2acykSIDxrV7rpI5gYOX666ozqlyLQ0fp+tc6IeHkhcyAmmJvrO1uCnWHheSqf//Nt376hU/Pez9LyR8ZZpQ/n9/YuJ3n8XPzYmueudmfDe6soUwENAMEe/P26kCkM4NF9TMHDy54t1EEaPha1K4Ud8f1NmYaytKinUVd/h9eu/7nH3yw6/YO788cP/4vL1/JJUwlAmu1cqXNh5np6WarlhdbzaSMtfcwFZ0B/ual9184cnh5f5McNkNUEwzdR4VcZaT6CTm2n0hC+BHj1ZXVVz6I/HmyQc1GvkD1cePjHavNw1lHgGqoWU0oz9BjE4cRja8jsWrkqakj9/DDDz31xBNPP/E4Aa6srr7x5jtnzp67dv0G+6TTmwsiAMDMnTS10pBZyvszkpoGLpiZmYmJEE2tP8gR0Tkn4ppeUt77EEKQ4J137Ji9qqiqATAzIYmpqqoZM4HVWR+IiOLDner1NuUX3xBAQuj3t1UNlAyiO8f0GTM0QAAGcIAeKUH2QB6RwdDAFFSjNjuuhiGFanoVG/2GgAhMSIxM6Jh8wol33rMnYkLn2TtOHJtIdItSVQPVEIJkIQy6c/NpZ2Fze1CQEzUgXXS99e3tX/7tvbu3RYsWLVq0+DigJaBbtGjRosUnAD/63/zK//c3//2YfC63cH31zoG5BRbtD1Y9mWPMBv2iKLxzRKVnBRKaATGnjpNO2hGJy9dF1SXeJ0kU0aIhqZKKiqppEFVTZNftzouiGViZu0g7SaoKiJybsBVpkj794BIAqF16/9bmylYmjfXFdeRWy78MVCQUBQD2XM85jyiqCmZEHMkGNUOEGD9gzMBXvjqraggBqeSIRURUSlEaxM1YqavMKm01E8U3/9gszrFIUjHXYNV7cpkLkdixizphAOCyJcFM09R7x/3+IMsLDYWKlO/T1erp8lJnETXD8M284i/Hz2pumaCykYgMNVq5IhERR65GDaPIzMxiJsdK5V1SzIg09OKo2EGrfQ7G2If96Rlx2ocpJawMBv/r62/8teefm5vBAfkjw+eXZvPfuDXGso0J3WciMuOJhdqbq7c/u7S3owgjfm5p6XevXI0nNryVPyAR2tB1TnRfJvKH169/efn4nqXMefen7z/225evTJbfUI42qtoPqlatvw84vmeiEcTsH757+q+/8Kn9+4CPxTa9kT96FXQu2vhtkuUHP7MC+sPAyiD7h+9OWlTfBXD8c7w1jY6ikXtjuaMeHaNdXt7ZKmZ5F0ekaaiSuxqWa4Oq5wLzkYP3LS/f/+STTx47dnRQFFcuX3n//cuXLl1e39wk53yaAgCLaMz1GhcclYtZqpANHcT8ByU5DITeewAon2VVXoFyNxEZA6ICQCSyq8U+ampgUJK/UatczgXGXYho5cOqnA82tRBEQmEqoBqJZ4Py+TFs3OqBgAAOKUVOiVNwCTIDQbXgxswQCEzVyttT+RRCQwPH5Bx5x4jmmDyT88xMjoliimMiQVQDLSQEyQk0BNBAiEzIhKaFgShCrzPXL0IBLg+QY5agS9n98u+/P3uftmjRokWLFt9dfIxeflq0aNGiRYtd8MN/45d+63/8Dw4+dG310tLq1vb2IJ/3TjZXjh1aTB1vbW2KmmO3uLjovTeAIkh8LfXOs3PxndZM86LwkMwxq2pRFNkgJzNnFkLI87zIg6Gxc2mSipgqEFGQTELe682RERhmQQrQINuPHDvQ7fb6g8LsWpblW8ECYE0EI2CDOEFDVBHVPATtdDrMBAgSzAySxFOVQAkAAJG9Q8QgAQAIyTlnpiKOiCPJoFoZZSLWBHTkqQFK0rp24agNl4kiCQ+IKCKqSlRJtZCIXJIkIQQRISbH7IizLDOTNE2Yib23ze1i0GC4iUyl4ag5vISpnRhXGpfHNmiTceYES+tnq1ZwN8FMRiQisXGIqRQLKlYyaC1jM0PFOiMiIplqTTTHnqqY8KbetOETvTeGjNwENzfh1gsAAJc2N//2a69/fDjoUwsLR7vdWY58dWVlkn8c2zLalPHDSP69+viXV1ZmIaAB4AtHj1YENDQ56Cnp82ZDgwkbgVUj1wx+78qVHzz+wCw07g8uH//alasVG7XD8WWVOGNKuLGRY6MxN4Kv6fhhg1/c3Pydy5d/6MSJWSqKJU2sUBjpqdGL+IgF0KUFx0RfDaNLvnsK6K0i/Pybb22F8IFLGt4NAYa9iiMcNEDD3b6aMRu9c9K4ZX5NQOv++Gcoc8maOWJCUhUCZKb5+flHHjz53HNPH7v//iyEcxcuvvnW25cvXwmFOOe6c3PxxgsIIhofso07PFZmFBDX36gqGGo1szi8yCpLoZnFJ118uonEY5GImCiIaFwKE6HD4McvZ5iVQSVInmcSClCN+WnRpo34au0CAnrkDvmuSzwQG6KpicUJ4ypOQjRAqjhzAwAkY4dJ4tLEIYEj8p69Z+eIEVUliASRkkI3AVMwQRUyQTDv2DtGVPLk094g6EAloMsK8ynnFv73r9+TmY8WLVq0aNHiI8LH4s2nRYsWLVq0mAU/9F//4zN/8Oxnf+p3fvu/+0sDLWSAPddd3y5Yt/IiFHkBYM45Edne3kqSTpKkaZJubm8BYjToICJAICLHHMB84pO0AwBgFlQlhBACoCmYiuVZIUEAkJAUMRSFiZEiEjOaFAMGONhJvvf5JwDd9vb2jfV8K6giikR9FkM0s4zvqLVcSkKeDZjJe4/sAMCzq9/GRVVCAARAzPPczIgo0sqqSmQ1AW1WLfytEFvJSv7UmrtExKzmpkFNS6FZSe4AIjFzCEVRhBAKQHBEjqOOTesaU+8RDIlCnquqTbpt7AAkBhiSKg0DhzJmmBDwWcNUtbkiO9LJVDIUtaa5LAEJYwYqKPXhSEA1WYM01APWocFYMNM27n5xNX/XPG0q+xxxaXPzf3rl1b/yzNPHZmN+P1TMmBfx6vb2tX6/uQUr45GRq65NJ4buE7VvRnlYHAGvrazmqsleGeQA4KGF+WO97vXtfqMSgFk190NYY/ANA4Kh2UEz+JUse2Vl5TMzZH08mKZfPHb0m9evN4ocZxRhWPWMETf0oliaKkwy+9Dko4cDzr564dKnDh+ecV6hXGtRlg1Qedjb6BRKafjzkaNQqT839O9Q9eE+PKDvLbZC+Nuvv3F5a/tDqwEbjT+8vQOUvT52F23sHtkUG2rX+7RNuddVNaqZiYBKr9s9enTp+eeePbF8/OCBxavXrp+/eOmdM2e3BoM8SAihCGGQ5fF2WM1+jgQfI0es9fsABmpG8b4NNPbtUFEzI6Y4DkUEAYmcxRy0QeKkclMhDyU1Pz5QCUGpfMSKikoo2edyTMc8gM0wyyIIwAE6RAKkKp0iaIicNVU1sSPHzEyemYmIkBmZgRldzOOAYKBFnmWZmEnUcRtAERQMidAzOUIm6HhOfccRMhoTdOcW0rmeEK7184BUBFs4VGR9atnnFi1atGjxiUNLQLdo0aJFi08SHvlTb5z9+lOLD95cOXsoA7OckFPoF2SmYCa6tr4GAKbW7w+yrOi7QZRL5VlG5YthNIckAyNi55JyeTCCc955jw5VtSgCszNRABDhInAIhRZqIb4wGyMSCpL4A3PPnDxS9Puvnbt67U5/M6gimNXvp1q/+2PJD1iR5wAYXMHOMbuAAihmJqJRmAwhmJmEEFnkPCtwwpETonxsZBl+KYCrtxOXL8ga8xaaRT7BwKL/porUhtWERORUVUQAlCiqlccoDXTex5Ys8kJkZumfaaylfs23KsNgRZcPRdGGkRloSFLrYsxUZMi+TKNVENBqqw1rHldWVHk+1wcMKexGgfuQC9Yi30YMe5x/bXv7b7308n/05JOfOnxo9oo+OL52+cqtwaD+lRBnlCG/ujKZfnDIJJX6xtEROkJfjp8Kueqbq7dfOHJ4ltq/cPTor56/MDN7uytw9EtThTr2AQC+duXKLAQ0APzwieVv3bihutPVjla9z0hn2VMpMcsGL1T/0Xun/6tPPT97e42HXjP1kfRF3JXB/BCRy0RvjWI1y/Y44kPAla3tn3/z7eZX6YOhuoJhWtSSN46EqjW5/5J9nnLFd9tFUwhoRAJAAzURnyQLBxZPnlh++OGHHnv0UTC7eu36e2fOXHz/8q2bt4AZiABAVFRDpFpHwht7hGBjZ0wjG+dFcZyAjnllzTRes6gikJk0jqjS+tVXX88g4WiDIZiaiZiKmppq1EsP2edqyNcPawQgwOj77IEZ4sM8PlstPh9dtPsCcEzM5DjmQo5rkgzRTC1oEFFEAFPToBpMBUGjAwkTEZFjl3pOHTuGbuJS7yIB7QjT+Tno9G5vrAejTCyXAFvYmxtj3Vu0aNGiRYtPAFoCukWLFi1afJKACABv/4uf/QsbOHfQ1nOEtc0Nb9Bx6F0CGO7cudPtdg8fOrK+sbm1tVUUxfz8fJIkg34/ujPULGySJD7xjpPoj+y9d4l3iWd2yGQInbTjkBAsaFFooWoh16IfBoOBmiQd3soyLHIq5Kn7DxxaWMiKrAjX89uDYCiGYoSgCDhcdVzmEcMiL4o8mEqnN5d2e0UQFSlCiMkDgTDyxVgt5ZUiIKFLvEmZZw+JkNB0qDSLr80x0aKKRM6IuBRW1/kGJRQigojsmJljRQAQimAG8XU4arUalMRQSU1ESZJ00tR5j9vb/c1iJg2qmVWr1IdUBNd/hIzywnFLySNQlE43y9LYStjgMLAham5Sno1DhmXW1NpY+kGb+LAfWINubahsh23YDAUAEDAT/fk33/y+Y8f+4sOnPoK0hHfy/P8+feaVldUGxwJPHzy4MFvVL99anap0hmrjVEOMKJstLx7rH+WHV1ZWZiSgP7+09NULF3RUvLxfzhEbddc81S44u75xfmPj1MLCniUvdbvfd/ToN65dn5gxGWLIjM0W+Fg7TyidsT5sRGAaGxzhzPr671+9+m8+8MAMVeGY0HaovB6N4buCTKQOph5L1tjy9StXL2xu/nuPPnJyfv4jiMcAvnnt+i+fPZ+L7H30/goeHRj1zBxM829ucqz1V2Kyn/ZtBV6eRYQAqAYg2k3TBx988HOfe+HJJx9HgDfeePNffetb165d7w8y51OLw8Ox5qoqpR9UI96K8B2rAeuFL1YlXQQYmWeNJUnQOL8MSIZqEn2ZDKp1P+XkphnUjy1mgIYuPh6BZhJUy8VAUJpGG4CVXwAcpgiITw8G9MgpugTZQVwCYIjAxEzkHXnPTISIDowRmRgRiCA6aBUhV1UwMRVEQwQ0BTAiSBw755LEdzqdxCfeua7n1LF36AkcAaF5ptQ7TZI7/WwjNyFEhOA6g2zwD36vlT+3aNGiRYtPHloCukWLFi1afPLwZ//7f/4P/tu//CY/+b35HwsQIDhMTHM0680vgNnqndUQFAiSTqpgQQIymVikYqOKNi8KEWUuSQRmZsfsHToCQkTruo5nVhUgs5LWobTTcd6rCWBg7xcAEV1fuTcPX/riZ+47dPEPX37nxlq2MdCAwyXINWEWiQSzUnIVikCUdzqp956dK103wUTVwJgYANRUHAMgOxYSrTIEVpwymGmk1hVKgw5mrsVcMQRVjcSXc845B6WU2LDyZGYX7ThK700VI0J2FIIgAjNLEFGJ5BmCIWKn202SZHtzsyiKvftsfzzIeOqtISpOBjFevoIaYOSgK6Pr6BxaswxVmWYajxq2SynsxPHV13dFt1kloZt29vi2usZvXr/+2urqjz300BfvP+buji3aC4Xq71658usX38+ieLwR0vfMln5wNcsubW6MOGnYeDtV5gjV+vcRUWJjusCGffvaympQdTO4cBzupI8sLp5ZW2sOiX1bcFRVTwpmpxdl8PXLV//jp/YmoAHgzz304Ldv3cri3E/c1CDsh41u4GfwLK5OwmbMdQnNi4iZNMemY+Ix/++5C88dOnQoTfesrj69dk2BUXOVkbkUvKuvx90iV6mzhTb70Ia2IXhufeNvvfTKs4cOfWn5+BP3Hfjwgrm8tfVPzp5/587ah1D2cHqkMVMynEYbWe0Rx2vDpqXsouYcS/nQKRfB2DSZc6OaekqnPExDQUTeuUceffSxRx954qknEOG906cvXLx48eL7l6/dzLMQFEOWQ8ymVxHKw9UndemESNycgotzf8QUV/aYRmcLBABrfA8VEAyIG6+riDG7LAIilbbRFjvvpwAAIABJREFUofKJAtDGzNJw2gSBwARUzUouGyubmdJ5A+sjy58M6AAT4BQ5JWJAjr5aiI7JOyKE0jkEY3+YqqkKmMYwJATRwISOmb1zTI7JO2ZGZkoT573znimWSZQwOlI28MSeEQEdMbIrDLZDAKaQ2/n0gYOy8ZVvvb5DP7Zo0aJFixYfa7QEdIsWLVq0+ETiEi0/qe92kvW+dFFZwNLuHGviyEKRZ/2+T5OYDihIyFW6SQKIUrsjE6mqqVbeFIAIxERMAgaEzKRJ8MxBgk+c8y6IEnrv2HuvRoVIaUVBxEbk+ZnuA4a03e+/cebq+zc3twstwKQyeoCSAihfjOP7rkoo8twxeUTvPdY6ZRUzYC4JaHUeEZBIRCLZ7JjjXis10Br/j43DFTddkrBR2QUGiBxV1QYiIiIxPSMARAoboHwFF3HM5ByHIgBidNaOlI9z7JxzzMSMgMycDQbROlprSWBTy9zE2DLy6uM0TWhJBYyxb+XBlfoPIerKImdTqrQREdBQLcokKZLMBkAl5wxD2sag1LWhjfNsHx02i+IXT5/+FxcvfunE8p+6//4O897nzIatEL5x7drXLl9Zz/NJNj8h+vRsBiCvrqxO22w4FM9Okrqj9HRs3FHydCDy1p07zx+aKYbvPXr0zNqHQfztCAP441u3/p3soYMzcLgHkuTHHnrw/zl7DkeNikfLQwDo8X7//G627ZR2nkSMIRP5pffO/GfPPbPP6nYoc0Jt/dGgkJncBgzgtdXV11ZX7+91Pndk6TNLRx7o9e5hGBc3N3/n8tVv37j54dwgGsTxkHPGkQm0pgsK2sgp9WGNWYK4HWuD7JG4xy6itL9AhDg/ayrO8eLC/JEjS88/98ypUw8t3rd4/sKFd06fPnv23J07G1lWMDt0LCLxLktxWU2VDnek9Oh7VdWpMc+rAhHF+UJVVYmPSgQgwOGKGESk+KQDADCMWWcNIa4CIgIArIykEKopXFAoMxSYmYKqqZlU7LMZliN53MoEAQiAABOkBChFlxAn0aC6fLZgdNiIQcS/HtBMVdEUARAVQTH6dDlKHHvvk8Q7Zu85SZwjZELnyDlyTFEWjSaR8vZEHsETAhKnqSFvbG3loiZYaHE4X11JPlLLphYtWrRo0eIeoiWgW7Ro0aLFJxIvvvji1178AdzWo3du3D62nCRubq4z1zskxUClAD0AACHIYJBlW5uqMp8krGpgg2yAiGknzYtCRSsCEwDATCVoXhQGQEyWCSGKyPz8HCH3t/qEuXbUO6emeZ4hMSKoBGBHLu0RPLF8+L77vkDwR3l27upqpmZSK8rKVfPY5I9UxYpsU0K315t3jhCJCBCdcilrrJlWQiKIhLmqOOcqArp+Va+UX433abPK61lVTU0tshiqoCpxL1ZMLhISsapEnXiEqgEYIjIzE3tm1dK0Mwa2uLiQDQZra+sb62uDOknd0Mm0WkJeqrOx9nkGgFLCGSljgEgrxK1U2UNb5atbnYjIXJIHaAAU8wpipc21SlxM7MwUEJEJ1EyNSiIeALRir6tQzBArDvqD2g0MWeyd+eyRPfGXO3n+K2fP/er5C88fOvTZpSPPHDyY3i0TvVWEt+/c+eNbN19fuS1jviCAUPnBvHDkSDJbFS/fWhmqK7EWe2OjXKytISpvhJoTq2YRqp4sTzQAgFdurcxIQH/myOGvnDkbVGsie79k6IhjgU3fNbZRwX736tW/eOrU5N4op8Th8IU/c/z4u2vrr66sjLiR4OgPgEOdGSTJ1Q+sUv81fUxG2nks9iFfCQDw5p3b37px43tnyzM53kHY+JZWH5ruHx8NMtVm4sF6UE2O53jEte3Br1289OsXLz0w1/vU4cOPLS4+vLhw15M6t7PslZXVb9+4eX5z417nYMTJD+X0WHPw1N+uEWn01LvUlIm8Rn81lz5MENCl3QXEhwyoLB448MTjj37+c5958MGHgsjLr7762tvvnLt0WRSAXDKXMLEBUp3GNuYQRPDO4WhayFpWHD9oFUT1ZENVES0fT4gU4xMzLDMTkIEpWHxgOWa1cmUAIiAag48lVldvIsEkZoUIIWgQNQkWcjDF+JgxAwMautiX96yYctADd5E75FL2DoAtirgRuOS0QwjUGHmgFsKAQL3jxGHiKPGukySdxHvHifPeOSJ0jI4pOnKoiRVBA3TSBEyLYmCE5F037TgCAgR2gG59u78lWigHKxJmkO2vf/3VyY5v0aJFixYtPhH4yGUMLVq0aNGixb3Dt//K57bvW5AekDvUS5PF3hyzIxnERe6iGgoZ5JmqddMumGkosmyAiIlPomhXVC1SqtXPIgQJoiqOOIqzut1OkiSDwQCQEp+knQ4xBRHnHROZFkCk5AbqCkpy6rxz8fpLb53/vT96/fpmvlGAAACRIUq5yniMCkEkSpJOt9vr9HrOOzCLsRERxryJpazMrMk8ASCVFFSEmSFxlFFXKjRkJuecVNR1rRSOr89aoVrSTVFMjTX/W9GXzMxMBBjTJDp28Y8IRhAJWZZng/6gPxhkmYZQOn4O+RKrSbPhnx5EULMq5YEY+Wmsz2zIa6Hm8BswHD1idGcldicrSfN6KqBaJt7IQFglsmr8vEtYHekkzbMTH41VHDUI8cTc3KMHDjw0P3+k0zncSReSZOrfbWq2XhSrg8HV7e3LW9vn1zcubm6Osc5TqhzlSA2AEAmAiDxhgpQ47jDPOz/n3bdv3pqa7xFqRS42tLmzXbaNHjLlPAQ08EQJs0MkxLUil526Zqw4G4YzUscsGOWOu849d/DgVghbRbEdZCAhV81FmhV6ojnnFpMkYTq9tr6/Kmy4oZpG+cDYVSddMdp7DPJmS+9hbF3Hj+N7R0d2NViGszyTgU5piYnWmnLi5HiuTyWkk3NzpxYXjnW7S93O0W73UJrStEsygK2iuNEfXNvevri5eXp97dp2v7qWD4l9bl4rjo+A6sa447k7bGhsrTP71bb+Vv5XfusQgBA4OhMx28L83NKRQ0899fjDD59aXj5+/er18+cvvP7mW7fW1jezXJHjnAsBAoCODqKGxflo7wzZ79Jpo5qjQ6xMos0Akag0nooeSqXMuU6hG/MQDM2xseHY0Zim0IqANg0qhRbBJIAKgiEMO7JewKEACIaAHilBToE7xB1mj8wGaIoIRqBUPkGqFMMIVLYvgjgy78gzeoeeMXUudY7QmMgRO89MSAgEQAhEyATMlCSOwFRD6qjjfbeTEiCSM5fc3t6+nReZQqEiBRVQ/MI33pna0y1atGjRosUnAi0B3aJFixYtPtn42os/gLxA3HEeEna9tNNzScoa1yCbgZWphiwaMYS8AAAmEhUJUoRCRFVE4j+qIhLyosjy+G5sZjEfk4ioGRJ2ez12Tg2SNHGO0AQQDSkPaC6lzlygzrsXr3/1t77xzuU7l+9kfVFBNKJCRBRGkiMBACAis/Ped3rzPe+dGWRZVoSCiIiZIgddLWuOYuQgoqoczWSHlKkhOSSK1HS1XpiZnVYEdGSmmTl6P+dFJkGkSkUYJY4xgWFslCpCjMkJ0SB6cTjn4vJnQitJAbWiKLY2t/IsC0VeceX1ZVYMLzUkmkNZ31Akh5GAHvsTpWLabXRjg7QdJUIMzLSU2SGBqaki1bS2wZCArjaADSm37wYBHeNoGLbWJ5UneqKec54oYXKIYpqrDkQ282KoMh6taJcY6uN3In/H2mDKn4ylarBR9+4E9OhhQ9n+FNF01SiTRU3F6DREHfzw8LEId8GuwU9aRe/Xh3qkosbVDvt7StD7Ldki47czazw7AT3RQROXD3sS0DBON08S0FO3AOzYs2MTH7DjeLY6+uaJCNBx3GFOiBMmNQimuchGUQS18R649+xzo2hs/jPhfT+dgJ7YsgcBHVHfPiP7XP1qiEBohADOYW+ue/Lk8Scef+yZZ59eXJwfDLJvfuObb7z+5uVr1ylJXbcrVqfuG7btEGaiagYwpRWrG21J4jZOqh5ARETkIBpPlU8rIkIz0OYTCsYGJgDUGQUBAUzEVM0UVEADaKik4CMEdB2agiGAA+ywT9GlyClxgsSAaIqqMXugUHkOxek6BGZkQkfoGSL1zARMwKie0BMhGCEykffMjGTgmL1z3rH3zEzM5Wqf1FHqOPEegMh1Ngf9m9vZpkmAUNyZo6T4e99stc8tWrRo0eKTjZaAbtGiRYsWn3j83s/9ZNGzpK9EtNDpHJhb4DxziTeAIoQk7bBzKqKqYEoAEiTLM+89syNENVXRIKGkmAGkCNlgAABgIKb97e3BYMBERQiDbJB2OoY4KHLnmIkQ1DnnnXcuBXRihEm3r3hjPf/9l09/643zF1e2toMqQm4mTVqofFlGAGZ27DyAAhIxG1jF3ZSeFYhIjI4dlkrqUipsQxYVzdAiq6RDOpWZ2bvIPpta5DhKjsbAQmEAGF+jx9ji+n2+FE1HzRdELlxUmSjx3sCIyDnPzISoIlubm5ubGyHPtU551/xzY+QzVoRz/J2ioK3BPw0xpHVHN0ZKYnxMxCxXZe0UF3APTQvqY8rf4gyFje/6QNiRg4aRjTaxZ3faEcd+qajq8eaatTicziGOUo1TyW2YUrNV9F5z2yRFuxNN/kH+LN2VJp61fBu/1nvAL+8SQ91cjXabqBHruZym8cgsgU09xoZeNrbTYXVFkx+mll95dsxU1NiJ9d7JLTBGz45OUUxWPXbiNM66cfub1lzj12iT9697Aqx+jA39Jit9F6TztFOG03sN9hkA0QwNTNEQDE2x1+kcOnzwsccefvKpJ06demiQDc6fv/DSSy9fv3ZzY2NTANl5ciwx4a0qqMYcAHVlBuU04wTBPPopct/Nm2B0agZAZCIGBDVTEcS4AAi1keGgWrxStSGVRUYCunRVijl2JZiKmaIZgAIqQEMmbYCAdawM4BB7nHbYeSAHxAAEaKqgWlLXBIBIAB7RETgC5zBh8kyewRMwGhEgGYIxgifqpon3zjsGUCZKnPeOvWPnOOacUDMRESnQlACYyCVdMbrTH2wjqFJ/3aMPVri//53vTHZ5ixYtWrRo8QlCS0C3aNGiRYs/Cfj1v/cTm4foobMBiFLqznc6qXfMwMwlq4DR0dSij3IIIWYQREConCjiMl8iUtWQF9HzoghFnuehCIi43d/e3Nzs9nrBdH1rI+aw11CAAROnSccUirxA58B3IFk8fW3j9fM3/+itc5dX1tcHRWYQSvthAGgS0IjERE5VEQmZnXfMXPKwhOUFUKkLjs6zkbYammQAgKGoqVWv6GAAGH08VCWucq7KKk+OVppWeU+rahQ6l7mVoiUnYbTmADCM7hwGQQITeecNDJHYRQI75lc0VckH/SLL8yKvyV+AHf7uqC04KjtuBBxzEYVmuw3br2YTbGxHSXAMKaXIR2ODF7HGeR8GAT0R1R7H3A0B3TjyLv+iw9GMeeOs6e6lTmNUJ7dMUtKTPO9M2uSZcW9UyR8wnhlKaMZpo67GTfG2WeUzUDVmzbruWT6MNn5TyTtCQO9Z2rRRNkJAj9LBU65xP1k+pxPQ0+Zt6v1NunlsPDcmTHCWdmsG/+G8K03eDEcJaLi3HHTz12iOBEQAoKqCgIlLep35Bx88eerUqUceOdWb64ZQvHfmzJmz58+dO5/1C1Fjn1S2TOVTx1Rx9Is2nCO0XdX1cVLVhmtfzDS6NiESUJnbIBpGISESVQrockCbDvu7Hl1oAFgmGAQAUxEJYGIWHx1WEtAwMiaimQYDMKIH6rkkJceAVGrE41oZi1kIY2oCRkwYPWPCmDhMHSUOHRojEFnlmAWe2TMnnl2UOYMxoec4a40IpqZiCkiiWoTcETrnfJIA+q1BnjHnQbe4n4Y563da9rlFixYtWvwJQJuEsEWLFi1a/EnA5iFavJWv9PLFfjcfbBuIwHwXXbeb9vv9oijSNCUmBAiqAJCmaczmF0QAhpLbSLi60vCYVBVz6vZ6zC5IcBsJIM0tzAeVAiRJEkLOB/08z4sQwHITybIBqKFLuBcePX7/oUNLg+1tCJJnawqm9QrkEZipiFpc8gtgROS9Y2JkIiYszSOwKAozS8otWDlX1+QQFkFEtdT5RQACgAgqKaohljaakXQlYjMLIvGNWCMXHT0rDBEhtgMhaUydpFamMxQ1HdaMAVXKRFKLi/MLiwt5mvS3t2UTtcjLXIxTtZENDEmLafLn6RgvZNgUscRaUmjNIyrmbUQS3cxJeG9Q8xyTvOYYPTlkUeoPE8fD6AeYIJumyol3rLr8xUbjGGMap9VmJZWPWJP4Uzk6Gzuv3LgbH32PcJfsMzTCmKGEaonAGF08awljLPkYT1r+iPLMscNsouPHiGYb6T+z8V4dA1ZfitnbbazGaihMCWy3a9zxwzDmsoApOv+RQTM8efp4bpw9U8+O3kbuPaounrI91oz1DOKOHHzzt7oDmiXUBzXbrsq6F2c1kMARLSzMLd+//JkXPv3EU08eWFy8cPHCq6+9/tLLr6zcvkPkDahMXSuios1i45NgpGIEBBqdVcPx2zRFo6Fh/s6oUy6LUTCI5llqCKCEFCcHq+QEzLWdtUGdrwAqXbRFJho0xqYA0Y+rOVVb3mERAAEr9hk9EMc1RDbk2cGU0KqUBYhgjsA7TBkTptRj6tAzMgChRdMsImamJEkSx2ZioHHBkBoGkSDB1CTkeV4UIbD3Chak6HQ7XedVrB+2C6VMtSfbar7vtv6P77wxOVZatGjRokWLTxw+pL+rWrRo0aJFi48av/6//Nn5LO2J75uEoAn5bpJaPuikSTdNE+8BVE0J8P9n7916JbmyM7F12XtH5jmnisUqksVmVbHZ7K7ulkeeBwMG7EfbsA3J0li2oV/gdwMDzNjCSA/9YkBvfrXnxQMYY9gjGJqBRxrLGEMyxh7JklottVpkF7ubRdaVLNaFVeeSmRF7reWHtSMy8nJOnSqyW2Jxf82ukxm5Y98iMiLj29/6VmBOKSJxzvnw8DAEjjEycZe7Rdsysz/SqioAUC/IypJz13VdR8wKkFW6LGJKQG3bLRYLaTswYyJGErV5J5T2MjX39ts/u/bhH/3Vj29+uni8kIwgJXeT63wJljxu0QITU0xxurMbUwqRXQUpYiL+oI7OC3sotKoycwgxpTSbz9vcIfijPfYvSLWkIUR0otWwPP+DqokqEYFZlkxIRGQ9PdDbT6OVvFDW0zPW0wdIhIToDYhIYE4pTZom53x0ePTk0cPFfAZo2Cd17P0xsJAjvbJ7ZL9BmwrogVJZoalXnWJx2GiFIQEABOrpCid1enm4rTANpR4vY7DO9Tw/nl7PSLW5JDRHVN0xO52uGG77bG3jmLpc23jMloEVW/Je68z6+DfmKgu4lXAeaNeVFk/4obrRs+c2aF6hL3G0ZcTcHWcu4QNaEzIPex3boo0OzFD/eMPIg/vkIZw0xvWTY73cmg30mKDDredEf4C2C5+XM9kroVeFzAabZ+xal8rnox3X+fa103Ktm5sK6OV36pjjuDK4lb8/pack3HiJy3/XljOQYHnJWu0dbJ4Z/QhHnyKhmYEqMQOC5q6Ifs2IMTbxyuXLX3/77Z/71s+99NLLXSfXfvjeB9ev37p9+8n+UdtlgxIc0y86jVpUAyhRMgAmooAISEhkYAqGgM7FqorqeFJtuNAPDDUAEKIZuoM0IjL1YwdQM1PzQ1l00wbgXlO+juiBN26XoWomptKT4960rp3KCMCIDBQAI1EAZMNIISDS8pAYgZFZDJxCiDEEwsiUAjIaoQVURmPEFNyDipidhGYiIgJVUckq2e96aB5cpKhKRBQ4hIAEBjrZm3JqjhbzDqIAZMBkeWqL/+4Pb510NlVUVFRUVHxxUBXQFRUVFRUvCH7xv/oXf/qbvzoXyZ0a5oNWjmaziNR1eTGbk1s4Ek6ahomPAJpJA4CaJZuBmhCJahFGOQuMBACIaKpgykWWHNRMAQMicxZTIk5Jm8lkfjRHsxgjGuScYTYTmaPmK+fPtm9fzNZNPrx/4/7+J/tzBBAEWT4OD9RqIUAlK4AxMxIQNz3PS8xsZiIyENAA4LYhzBQCxxSKJ2ZPFRT6mFiNzMzp5PKMP7TbkzJRA/QMBlFJftj3DVRBQZ2hLtJqK5OFiKioii4zV1NRQcQ0SZPdHUDIuTOzFYqrDNxwg4/cSqYuc2kNhYfMjOt1usDO+qIr9Jfz78fTwlsJ28+ClQq36RgH9CT4Nubr2bu1ztevf7Da8LPUv6zAxha7z9LDcYvjpm11+MfShXbMNP1MgaMXI4r9mSoYjvlow09naFuqNMNjUxE+9ZxY7fnafscVh+UKBML63mvf1ufHM57Pqz1b6cznjtE5M+KZe4Z8w596vB5i46m1kbnzej3LlnA4obSQtqYARkST6fTsS2cvvHL+W9/+5ptX3rxw/sLDB48+/PDW97//g08+eXB0NAdk4gTg64YAAMVaYvldLQt36On4AmDvf+yxPn55JkQwXnUzGV/CoV/CQSZSNRD16BtiBr//mqENZlNWVih8T5dFF+MnADADBV8rHSTVy3+XxwABCDAABaQAlJDYkMBcvO0LwSXNIGJATMwpcIwcCQNjICAEBCtzg6CAaAhqWQU6BcgAVkKePBdiobMBAAiBkZhjDDEERkIjIE6H8/kcUFA6gwDUYvjv//VPTjydKioqKioqvkj46/7pXlFRUVFR8bni97/zKwaKQIuubbPuMlgHs/1Pu8UsBd6dTs+cOaOqBwcHZ8+e3d3dTSllkZwzgKXUTKbTGCMxAYBbcLRt65G/KSVV7bpODbNaJ4JMQCgiIQRmbmdzVUPErm2l60zlcP9gvmh5uquTMweQ/uj71/7k3Zt/9t7HgpAR5uJ0t/tQ98KwgvIc3Eynk52dGEMIMcamaRpAWCwWbrDhimMRcVeNEII5yWBmvaX1eHIQ0fXdLigzA1dsMbOImAERikjOYqZE7Ammit+nSpbcdV0IIcWIhGBFJG5mnhcRzKhYduBisUDEGCMxd127//hxns+l60aut8telQ0DpbJNAU19scEMeoN9do5jqM3MFMxVhH2SqzI7PStRxNyFx1/W8/l4QG/2bZ1y7SPtl9TXVvptk03bKIYbVS0Z+w1l7cre/Zt1nelGV9fLrI5u0MVu7LhNBrv+YkW7aT1HBOt62NVhr+34VLHzCerX9RR2T69qK41/zNLBU+paezcQiKtK3ONp6bHV+dYWt/V21EFcTuhwyE7V4pZj7V+l9Qq2HKnRQdza6XIle+ppufrdGDd03Lnx1GN98nQ9O3D0dzi4uNJ2oTGXBPToGzO+NA0dc5+lDbp6dNlEAERUy6YCJmWmVAEsNukrb7z+9tff/va3v3X16lUO/MEHH/7JH3/33XeuPXlyGMKkmex2WRAwxqAqRBBCKKZLvXzZl0LbrvPbyqRpPHSmlc4AENnMVCXn7KE0J06RIUJgEtWcs6uEETEwExEADW5PHmWDPUDdhkpMfNHTB2ugAqbLBR3U8ZwSAhkEcL0zBaQITAaeo5gRmZAJCZHQUuAmhogYCJkRzQgtsCEiEbDnSCBCvwtm6URyFhFR6UCVAgdm10c73xyZI1OMflfngGSEC20XkueAyrTIFJmU8/9U2eeKioqKihcLlYCuqKioqHjR8Pvf+ZXctdZ1GVANJ2ABIM8PyIyJVJWIYoym/jCNIQQOIcTgz7QcAjETU4qJCHOWGEOI0VRdeGWIYtiqIRGgSc5mCkMaJaLcdabKRPPZrF20RsHSRNLk04Veu3H/D//iJ9c+/Pj2/f1DhQykS6JwxGD1phzMHFJqppPJdDqZ7rgcTEUGkwp1O+Yi2kLrzS6dggbPM+U+11gqLCHVqipmAIPPBhERc85ZcnafZzOLMToNnXMrIoAQOIQQevo7Q5Fmk7l+28xTSomImSFAahoiFMntbLaYzeazmYoUNd/Ygrl0saggNwnoYvWJS2YOl+WH+Vu1Pi18SZkT6IkTn+GiWV3hnfvefP4ENKysL/S03BqbNhrIstxW9tk2im1gNBPrO55U2gtto4lP/tG4Sto96w/Mk+hI20IHb/WSPqH6vnfHCn6fgpWZO56gHJp5rkZsfZJxy6xvXaHYinIgn3bgAJ53WjYJ6i2LFttI3vHZdRxvv75ms3paLolaWz11T+jcaXC66TodcO3vkoHuo1P6zT373G8r62PLK9Oq3hnhmOFtIaABDaC3pDAFtFdeeeXypUtvv/21y1cuX3z94qNPH928dfvdd6999PEnjz89EAHiGDiqqGeXVckIFplFVYoHdDkYap68F4gopgh+PUXwFUQ1UxGRjIS0SUDj2tEyBFNRcY+mMpzecMNvb+XepiMVtq+2ipkW02fPeWtDJYW4HuaEEANiAIxAETkgB8+9YECmgYEJAmEgJCJGi8wxBEbgEvsDxe/DSkIE/4umaCVPISIgGJoiaIycYpqkFDwbISEjBqYYYowxMINImE4P57NHXbtAyIDT7mwLi3/03R9sO6kqKioqKiq+wKgWHBUVFRUVLxr+ve/80//zv/4Ps5qIcAhq2DRxGl+ybqGiR0eHyJwm01k7W7StiKSYUpMQJiLSth15BsLAKaUQGAwlxdDlnDMhhhCBUJGNGA0QkBBVTUWIkAgBDAKBETFNcZpiUrAMprB4+bULezvTaQyTGAnu3nz45EigG3w3YJNSMMlZVQGBiJhDnxjJ/DkXAN1VEvoncSQC7NlWAwBwkfTAZYgYke+4jGp2Fp6IILuTs5pqlrIjsxJiV2TRpGhZFAu1rQCeuQk9OtsUREQ0A4BnSAREF3vRzo7rr9vFInftFhbPxq90/VNAGxsE4ygkfbzjKgM94pTLP2grOxzTgxOo2ufGRp3HNoIDwXQiGYbH8VDb3v40KPXNzmxr/5nrOb7mHqcYzOcy6m1NnySP/UynzSb1ab2w/TmbOzUeFleWAAAgAElEQVSdepIXxzPi2Q/+cXtsHMGTh/vZeeOfBvv8TM0DQu8b1NOnGwMuJv7H1GCr0zVawqLAMaadvZ23v/a1b169evnypcl0cnR4eO3aez+89t7712+IEVJkYgXoRBAATS2rqqCZSlZRFVk21i8ymIEpmhVPqeLUgai+FmkKhiKj6zka9AuKo8qcyV2P2nH2mZCQsBfYl2LLNcSBd1YF02INXaYUxicNITBAQEzICSiAs89EgIRGyIEssAWyQMTkRhkUCNwV2r+MCiaqoiqm4v8XITB2lXTgwBQYmSwwpMBNik3TxBCYAEwJMRCFGFIMIUQx6Drt1ASolRx3tcPD1O5uP8IVFRUVFRVfZFQFdEVFRUXFi4n//e/++/vx5T3dnzBNQtgJiTRb16p2plqedtUULOcMALu7u12X57MZufaJCBCYOKUmS5acB+0wAFFMcWfX1cGuJyY09uRLJggkal3uyIiJOPDh0cGT/X1spmHnXNh77S/fv/vHP/jJv/zD7330ZH6YsQQJL50oeupFrejYCEOMoZmkJiFh1+XyDK4AxTm0kBb+4Fv2GVkk+2DN1HkmFS2qtJ7SDiEAQBZxQTR4sPMydVTRvHkNSH2OQ8Ccs5lRaRQJKUuXc4dYlNUllyPjzs7OtGkY6eBg//Hjx9J2rhlfUegu5Y7rKLoyGP14QVqX+RY/6rLFwACMwM2ye7bdbKm89Pqw10PrILr86emgAfpxrvLnW8Sj/QvYzFK4WewUOmXbWtVx9fb7lJPwtON6WsEVH4x14ffTOv9cv1u32mU8c1XlIJ1mt+fp6gm89nNTw89qJXH6htZ1zcPqDqyf0+s61zUp9Cl6OHxZ1lvctuuWs+vpJ+QznOGnxrbatqworTpBn1DD8qJ3TFfHF6v+6CChoYEp5G737N6rF1+9evXq1W9cvXzpkqpev/7+n//5927evP3o8ZNOAUMDFNysCA1jjGAmXQZQUzU38R+vC3qDhEQMgGrmVhtmWOKBkDzixsNpljuh37c2llvG+WAHkw1/RcN9ydRARVTEtKQfNMugNtI+a8++67irCBAAIlKDnChE4gDIgEX+jMgEDJlQGSEwMxMTBfKbWyHTPY1gVvEsviXZoHPKCAExMgVCJmgipUSBMQSKgQMHRDATQghEKcaYmtBM9g+Onhwunph1llszJA2N/qM/+GDLIa6oqKioqPiCoxLQFRUVFRUvLP6Hf/Bf3k1X/p3DPyTiSeC96YRVGLJJJ132x+as1nWdqU2nOyJ5sVgAgqh4oj9EMrOcs6rGGERksVjE1CAHAQwhxBhCCERIZOV5lEnVACmE4LmUmhTbdjGfHQFHiDvYnHmS+frHn/4/33vnz67dfO/W/Q5AkAwJXM411kMPMf3MFGKaNBwC9BI5LQT0iJjpH9hdTQYAxMTEOfdscolhBiJ0y04v6dy6mg4cW08HFDYWoXco9WBoK+NVU+u1yMTcxARgqiK9CbVbVE+a1KTGReU55/lsfvD4yWIxLxy0j2eT/hqRFO4iaqUHw6cbKuA1xmuVMsSRJtpnY1DJWd8BHJR1Q8d+WrDTy3S3qj/XyL1T/K5bIfBHXHu/caNDp6t23KVn3aM0cwpu99lZ4+MpTjd0Gd6VTqwWWXbutD1cNrsynycV9H+eUu7EWd1+Ej2fkfFn0kGvTWfpxjYu/hnY/LLDFvL2uKLHO31vdmNdMPw5YBAeb1S78h1euWKvbFxO41YW+7h+msuIh8UBlyYDwu7O9MKFl9+49MblK5e/+uZXQ4jz+fzmzZs3bty8devm0dG8y2ocFEnBM+4CAnFgNDCR/p4hw9WyrPINgmdfgzUtnHdZDVUoi5BUQmH6IRsagG3LHzvkNSyy514P7a4WSO63YaqSXYRcbpiawX05TFcO6sjcHAEIIAEl5IZCIg6EpMAAZIZQUg4G9swOwERMSAhUvhSGHoFTvECAiAiJ2X2qncgGRggEgZAQImNkAFBmDIH9hkuMgSkypxDCzu6ik/v7s7lpq5AzAIqA/eP/78fHHOKKioqKioovNqoFR0VFRUXFC4u76co3Fj/KHEDB1Di3L+3sNqwonebMFAxQ1HInppZiMrOmmXS57XLXdR1zMLP5fG5mLr7KOc/nc0DUrj2azYkwcIgpuTEkmIUYUmpyzszhzJmzWVTUctMQWqQAQO18fvDkaOf8xbdfP69/+5uLhTx+fPRgtpiLKSB4UiXrfTZxYFgNVFVy1xIApCZ5mDMiA+DygbuXGyNi7rrs4dLWW2OYeqokAAhFtgVqoFjy9SEiM0kuWQ1x6EGhZA17RgEQJJdYbA5FLg2ITBgCuWd0l7PknEUMIDBP0gQRJQsYhBDPnkm5zaqWc1e03EsueISBTMIl49Fv6V+sCC/XgO414vJp14rDYE+ybM2cD1mSsSuR7PhT46BxIHQ2uc+tdLOtvt34/FQtrkzYuNIxD7bJlJ0OxTWiaF9Prag9dedPVwD79YWTqz2hwg155rPNQ1/zeHFkU5B7ah629+I4YcFiZSzPnUbvmbw41qneY6Zzvdgzs8/gX+TTlz4VB/15Gm4MOJ59Pk4TvaJo7ndfDuDUVLqXLtc1A2BEYMTUpNdee+XqN69+7a23Ll58fWd35+aNWz+8du3dd959/PgJAHGIzSQYUSfaifjyHhECGqCrmx0RQMEMzSNdhu71d4lyLfO4l43OWb8og05Abx+ZE8zg13tCcUtooH4/v5EN54KZCahAIcdhm3FT6SYZBoCInDBE5IDIBp6SEQCQCsntuudiKIUltwNKWSAmREIMTEzsltDM7BkLUY3ACIDJCIE9XUNWAwVFt+TiwBSiIRiBMc679tHB7AioE7BmThA18z/+4x+e7ohXVFRUVFR88VAV0BUVFRUVLzL++a/9J6gaVKRJKfCre3tn9naSSsPYtYssAhA8Y5A/h5rZ/uETA5tOm9lstli0ZsbMiDCfL1QFANwmWdREsqqWSGEE/xSRVBWRYmo6UTWIMZIZqCCSIiuGBXBHsQvN3U8XP7714F/92Q9u3d8/zKAIAiBLF8xCTjgZoAhIzCGElEKMKaXJdIeIi6bXCtNKiDGEnCV3nagSAhF1nQAYM7tPdAwRicBQTSXnLJmQ3FlDRFQEEZnZy/eWm0XR7FYknmMQ0HzsAODEleQ8WH9YbwONANS7TnvNRBQ5dF13eHi4mM26ru25gG2h9S5/c702AHiirSUBvZqha7nXkvkYYtJ7omapjOs/NVgmKsQ+z9XPQAQ9tLIc+FaXjFGPt9Dtz0ilrQxnjdQcGZg8/6/EFSXnmIHFtVKnoYlXa34KEVl6f8o6T6xteQie7/ifIFseVfg5jn2o/LP+vC8Nbfsu+vaeS1z/ZgzfyBO2QNn1OXs1JpdXKPnxRRNGyQmHwp9HH57ax9W//Z8tbPKK+cYxx/U0a0zLbxciBKTioIGQUtzb3fv6N95+662vXnnzStM0h4dHP/rRj6+/f/32rTuz+RwMA3MWMyKIMauKCqghEjKx88ijnhEhIZiqh8WoKsCYoe611/563MchumTZa8Rtg/HkuWV6XHi8krrVzBTEQEVN1K2fQUBlud6z3jYgAgFGpATcADn1zM5qmwbEwFQSEbuYuSy6KoCZKaEFAETzFL9FEw3GrpIOFJj8N4SbjxAYoSFADJgCpSaGwCFwjIFjwBBElJgjx8ez+UG2TvCQY4CWwqI6b1RUVFRUvNioCuiKioqKihcZv/Sbv/N7f+8/shgY0ZA+nS04NGFvR6U1QEYOMSGSE9CuslNQQGuaZAb+dO2p84hI1RBRRTyzkpmpate5OSbk3DnBms1UtW27wtGCgYpJJmIgVuB51hYYm52Xp803Lr28/+Ry4o9+cvtha9D2Iq7hedof6ktGPRXJpV0AiCm5PSYgmoFaYSKd8CUi9IxQhN5dIrTydG9kPQdCnj8Jyf+vKERIyEwhsLdFaqJg5oyDy4lhSTQjgIELn91qGgyICQCKVbSZivrklPhlpBBCCMzMsxDm81m7WKjknvldhWuW1UO8cck7nUzHbcqpFcYUBXpVtiSgj9//GcS8z47RiErDq4rI9cLreHameFUtu63Gz4gt1OUmzQ7wHNzu55gu79QtPu+OSzH4cRU+o7r8FGP/7OxzaWhTwV0+g+3by45P3/LczO8wfFtNzjhmn8ctHseff5Y+PAvG3+iT29vUxm++PUWXDQzUTJlpd2/n4sXXrly+8uZX3zx//nxK6d69e7du3r527b179z45eHJAHIg4m4qbD6GoGzcbABm4ddIai4ygWFyaB3smxY20hBuvy2V2ZSzblgwBwJMWegmkjTLus2FQsg4qgK4ce1x/hwBkGIgiYgAICAEgIJLfIhEJkZmIGYkUUYelXFMwVVVGCNDzzmSMQAAE6muq7g4NjEwYCBmAmZiACFKglELTpBDYF32BMJtRiGJ4eDibAc4NLOSk0GL6n//g2tMOcEVFRUVFxRcbVQFdUVFRUfHi4/d+45fdSEGAdkJ8+czuDhHLIhLuTHedvwsQDEDNgP0xXhaL1vMTOoUqKjmLqjKRAWTTFCMAHBweuBy4azsAYObZbNblbEjOBhuiSKvShhDUsMvWKbQKcwFKO5B2jjJ9769u/N9/9FePRQ/U5utP1dA/Sg+P14jMnNLO3m7TNCEEZAYwVTUxNGQiVRVRjxEmoq7rnLNWEc8Z6BaWiKhmRccNgIgiIipIxIE5BNVe/6zaW5GYqokIkftcq5mpWoyRmIpOGqzno22Z0tAMzHwvZgY1ZkopLRaLo6OjJ0/228VccltsTMcqxzIHWFTPxKv6wWPoDBt8fksOwp476wnbQcCpI87fP1jzA1nTTVdUVFQsgRvvVteQNkn8dYuQEkWyvcJtG4aKRhpvBRMCm0ybS29e+ls//2/8mz//85NmMp8v7t//5C/+4i9/8uOfPHr0qaohMhGbQhbhEIBIAMvaISIyI5NlWRr0g18qtXS9X340UxNZ7dKQEXe1n6cloA3MKyQA3vi4d8wwKUS4LxmvOW/0C7EEQAABMREzICMkwoSckLkYMi/XUBVRDKy4YJmpghqoERibMhIjBgIiCAQRITJExhRCZIwBJ4mbQJEwRvL/UuQYKISIiGZAHLPq0XxmnPaP5odKGTm2rSTSAP/jv6q+zxUVFRUVLz4qAV1RUVFR8aXA7/3GL4uRARMYGJylINJRd3ThpTMpBELsOkV0l0YiQqQi6RXJ4ImWiEQk565pJoi4yJ31VKmZqcpivnAmV0SySNsJEAGSmEpus7QxRAXosoiCKAiwICtGTLv399vrdx79wZ++897tTw4UMoCMH+HRn6aHB/tCE4QY06RpJpMYIxEZGEiRqImIGaQUmRkAc85mRlg8oIld+4VmWqhqLMiSVdVTLHkORigMLlifeBAQVBQAiEoBZvKchd5f69HvawBObSv2s2mihNiHPjMiHh7sHxzsd22rIksOek2IjAgU1qPrj6Ezej6npz/GBPQyct0K3VzSLRZd9IqQ8mfkxVFRUfGFw/gqNGzAbQX6P1sU0dvKH7+hh0vBi+kFETYpXHz9tStXLr/11puvvHphd3fn7p2Pbt26/eEHHz64/+Bg/0ABTNEAiYMZqAgiG2IvbTZkosDMrFLS2A5tFaeqIX1nWWpc8dvefiHectnEDQq+lOxvIuhmVp46F4uw30xFpesDhJyA7vnm8axYYZ8jUkKKRDFwDMyAATB4KI6BiRZvKQAXVPehUIBgBIBWFNORKTK7i0YkjGiRIAZMkWPkFGiSYgoUCELgECgyckAmKH4lgFkhGx617aztFkgZaW4dh8X0cPIPv/v+cQe4oqKioqLiRUIloCsqKioqviz4nV//z81UVM0UO2CVncgXdhObmEgWc2rUQDlwamLTNETYtq3bFocQRaTruul0Ssyi4vroZjLxgOWcswEQogGoattlNVADBcjSSVFAW5c7d0VW4E40G8bJrlDa7+Bf/uu//LNrNz64/+n+Is/FBMjA1ABKMHKhRpd8KFFIKTVNTIkDM5EruFQ1i5hZjNG5XRFVVeq5AzdV7qlzVSlO1oQoqmpaMu8VsfCSYekB6n4frphDZGYRcf7dy6sWL+ve/7R4ZyMUpsZUEZAZm2YyaZpmMlnMZ7Ojo8Vi3i7arm37zISwwkS7AnqdgKahh+MjPnpjyxSDw2c40M5LArooq/so837vSkBXVFRsYo19XnF2Xi14IsV8wkfr6mpPpFpY1/LGbGdneubsmfPnz331rTevXLny2quvzBfze/fuvf/++zdv3v74o481CyKGmMzIDLGPUAEncT0/LQIQetRMWbOzPoLEjZuWa6BldXHo2GAjMjDiS9jW6yatbLYSkqI2XHjRjZu8Bv/PNKt0UFh8v6aPIlpg0D4jAwTARJyQA1NkCkxggGakhoBgoFltrW8IgEAEbqlBiAEwIkamFCjG0ESKjBEtBoyBUgpObTcpRSZEX6NFJr+Fatu2qgpAyiEDfXrwpMOYCdus8tZP6Mm5//X3Pj32XKioqKioqHixUAnoioqKioovEf7Zr/0dMzAkldwgvLI3feXMS4eP788P90NoVK3rusOjQ2Y6e3YvxggAi8WcyHP/BVXNOccYU0pp0uScEXE6nbriOKUUU3Se2tQQab5o2y5jYDURFWYSzYvFIsZEGCRrm3MnoogQGwg7dz6d/cWPbvz+H33vxidH9w9zxtCZZTNAAhukxGOTSyqkcAgxxaZpoNesiWgWMdUQQowpZxFVD6k2M5HOgJCC+yC7yoxc3QxQRGEipgIw6K8BCYnZVE0NmcDENAMxIhGhSjY1KGHNOMifp9MpM2UR9wAJIRSWwclkRERi5pRSk2IMQUX2D/Y/ffSpdJ1pBrDiuaFa+B0j33M0D73w7pjcVogrBLQNQfCFROlndWkrO9Zur2zc8rqiouLLiOPY5+HPmv/GU83Ln6Z9NnPfCJVsCOjXQBWT7spbX337629/61tXL1y4sDPdWbTdO++886d/8icPHz5ctB1zZCYiKg7GQL5oV5hlQuSyhqel3+gBQOreS71JEfbu+divK9qIovaXm87Nm/yzVzkOlAEzQoLe/sK1z+NW1NQkgylYr8WG3sJ/fCsothsUkCJiopAoBCQALX7Xoqbq9w8zv+sxEwf3pDJhNGZIgWLgSBAQGIHBImOM3ESOEQJriuy/BJgDM6fYIJGIx/kogKloznk2OxJRIBbihZrGKAja8f/yvWv/7t/evfytw9/6raecExUVFRUVFS8MKgFdUVFRUfHlwm//2q+IiqJFxZ3Ir+7tgMHRo0+6rpukNJ00Bwf7OXcheJ5eT/eHAJZzJuKUUs6ZiNKk8YdnIlQ1Mw0xhBCZg6kyc0oTURWFEIOaqmkI7ukhnWQADCF1OXddBkbDIBhmFj5+dPTezXt/+s4H73x47/5Rnot21it8V/nQIkpzhTIREYXATTMJMQ6P9YjIxIScc/ZgZiYCxC5nA2eUiXoyAYeEgWai4lHMS5nZIEZ2Ew8iAANTQDQAM+31Z4BIzOR1qlrTpBACErm8rdhrAsQYzaxtFyEE9y2JgWOIMQYRbdvF0eHh7OhoPp/7UJaDNuyzEUKZlhEBXQLg16PgDcF6xnmNxR+MOQYOeuQWvdV8YyxCr6io+BuE4x5tPr8v7HYt8zr7DBvs8wk1PnVbsSo2K5SsZAAjRo7h5ZfPfeUrF9/62tfeeOON8+dfPjo6evjw4e1bd2/evHX79u2sYgaAjAgIREhmnvkTDcD8eo59UkcD7a+jiNSrq0u+QSxXUQQb7gZITH2eALfsMMLRtdpfma2t2BmgAZZVVZV+jAQwrLSamnHxiTI1MRVQ98kYRNbr9aLz64gNhYhEBgzIg3eVj8L5agMEJEAmZubAHJgYMaAGtEAQAkWmSBgZI2EMmAKnyCFgCBCD22shIqo5kR3AUMzaruu6TrKYeCwRpZ1dRDzKXQ6cEbMYf+P6rXfP/OEP9o8/JSoqKioqKl5AhL/uDlRUVFRUVPxM8Z/95j/9J//NL7EagCwE7h8cTJhpspvzY2Bqpo2ZLBbzruvcRpmIzFRE5vNZCJGI5vOZqvFi7s/GXdcOz8BERMRmyhSayQSRkNi5bDUNIbjE+GgxV7PpdCdn6XJGIjHoxICbszH9rbcu7+/PDo7m7d1HOjcxM9t4pB/+ummEqqq2OccQMSYiQiImImZCAkCXb3sPETEZuBzaPZ25yN+KctlURQQR+0BsM/XEjAB9EioiwsK5uIu0eM2qy8yHLgxn5hBCjBEQTK3rOqdRmqZxsVhKEQBcO4YAHCil2EwaDoE4AFHuOhHRolS2VQLIp8GWBHXPTOBqsSFCfG3P/sX6DG8vVVFR8TcXJ5O8n/vX+PTs82kqOWmbc6bDQiAThsCTSdo9e+bNr1759s99+7VXX5tMp7Oj2e07d65fv379+o2D/UMVCSkCYs5++RdCUHMWFwYCuoSAuOtQWYtcNj1QvIPuuJDEZn1MjKnq4JIBSOtrfGuLgcUEipxTB+19Nmh0bUdAxHLzMTXVgacelgw3myBwxhkDIrtRlJqY+2AheaslSMdF4BSIAhGzv7BIHMkCAjMFxkAQmZpQMgrGgEhA5OuvKqoeaSRZXZatAL6oLJ2gKhOlM2fMcJGzhtRmQSKaHurDc5d/7lP4wVPOjIqKioqKihcMVQFdUVFRUfFlxG///V8AQg0QMjZAZ3fTJKRgi4RAyCJ5Pl+IiJm51FdVuy67NCvnEmeLgQCsbVtP6Ne2LYAR82KxyF1WVURiZOZoZqrGgRAZENWJ7RhUvTZTNVVbtBlCMzlz7tFcP7z3+I/f/ckHDw4+ORJFMgB12qB/8jYoYt/BuBgAUpo0zXQymaaUQogAQEXlTOajyNnMOAY1zTKw0ACFV0YzMDVVGSTRgOiCOATwCRm2InlhFRVPW6ilQkTEnHPbtt6xwlkjuk80EWnhHSzEiIgqJQsUQGEfmmbCRCpysH9weHgwPzrSpdgZ100weofonghC6+PicanIs+L83Mv9NpTQYy8Os3EBG1gP2NiloqLiZ4OnPbmc8Pnm+t0zNXqcvfwK+7xqBrEqzwVYVU+vR2mcCDX0hLcIiMCMF155+dKli199681Lly69/vobBweHH3388bX3fnTnzt0HDx4uFi0hx5jUVLJ0uQM1M0Akg3WTjP5WAivrdGP//XIFVQ95Qb9AE4KaiTsjERIiESKoqIG5mYfDFcZ9A0tDDnLDJFMd5R4cT6/mbDn32mfp42+2ENAIQAhOPbv2GXtOm8olv7DPXoABGZEBmMn/IwJCcItnAiBGImS0xJQCERqYqYqaEFmKjL7J0yKqBmZXcPvSb+QQwCIzpebJop0ZzRFa6B7td6+f2fut7/34tMe9oqKioqLiBUIloCsqKioqvqT43379FykDqIXIienVM2d2JlNYHDKA5+ZzlZc/wLuw1z2gidkMOsmAoKZt27o2rWtbM0Oitm0li4GpGBgwcc6SsxAhIKqhqBkCMQORKsxmMwSKIeYuKxDGxtL0QOjGg8d/9eG9d29+8nDWzXNJ6rf68N1bcPTEAVGIMU0mu5NJk1JysgCLubN5/9WMY7DeWLM8/Zt5PLXXOM4fWAiHsl2dbXdBXVFMl5R90Het5IvKIrnr3Eu0y93QE++UiLiGjpkBUEU8o1bOGRDcFTowMxIASs4H+/vzxbzrOigJqEYYvcU+0WJvEo1rgj6ENUH5Uk2+WpeNHKJHn67RWJWDrqj42eF5Cej17+jpv7NbtczHaZ9x5fPlxWHYjutlTgUDUTBDxMnOZO/smVdfvXDp8lcuX3795fMvM/FsNr9x49bNm7dv37l7eHS0aDtVI0RGLquV6rn9zLSoj1cGg4hEqypl6G36/Xrvnke6HM4wQDUAKl7+/RLjMl1BYd2pt9coO2GpohRzFBraO2kGZipiIqAKoCXMZfUeOEw6ATAiI0akgARSxNzUU/7kKQyQAlJCCoiMQKbsW9lHYIHAZ4IICYHAUuAUuDe/NkQgopiI/NZaVmCVey8rQmKmyDHFSESzRXdgNlM7aPF3373+rdfPXvvoyekPfEVFRUVFxYuEasFRUVFRUfElxX/x3/7ub//9XyAiVcpo+/M5ETVxatoxWArMSAbW5bZrW1VtmkbV2jZPphNkziqqKjnnnEXVuV1/ZhcRAGDmruskZzTosnRth4iiltW6LosZMYfo8dFdoLC7swdgXdcdztrAeubs3huXXt/ZmYosrt198uCgXYjJyghWuQwDMFDJnQGA548y53YHIV7/mA9Z1R+XFUBURcSZiRC4FzgPlYLqkiMwc7m15ZxtxOwSoYiqFQNQVfU5MbOECABd59kWsUkREM3AZ8ml0maWu0yBiKBdtEQUUpzPF4QYOLx87tz0zFkkwn0yPdSeq1iZiaVS2Va3GCCOA8ttfa/+D6INFh7uNOLB4s53r1t8WNlxLGN8follRUXFabDmmXP850/BKtu66epz0l6jPqyxz0M1fUBGeb2sf8T8Wu+scWxjOORHRTQiCCGcP3/ujcuXrl79+huXvnL+wkvtYnHn7t1rP/zRj370k3v3PhGxkFIIUbJIFpEFMhMzhwCAqiZZihdF6S8CABJR4GGR0VfZ0BSgyJrJE/T5pbDPOliyDAAVw/2SURZLhlkAd5kGAI/v8Rat8MVIiCqiVsTTagaSTdVErXhuKJiB9j7Px3ioUM8+B0DnlwMSoEK55pfbJCEyon8aiCICgYEpImBvDI0AIqpiAMCEjGAI2ZgsIKJncYwhhMDEw0KqRzep24cQFRNqIsgq7Ww+R5wZzBe2e+3mv31m908q+1xRUVFR8SVGVUBXVFRUVHyp8c9+7e8QKaFSDBMML+/u7e3shjxHaT0vk6n487B5CLJBSCnEyCH25o/qD6Nd13naITd6NtMsuain0b2hLYu22Tp6wMUAACAASURBVGlkEzViQqRF2yICUwAEEVksMqYEIQnxo8PFrQePv/vu9b/88P57Hx3kPrDZioptTHiYO0wgIGIgdn47xRiY2W2anfPtlWmIbuo5onOLqMuBiISqigAEpKqqUqbAwEzNdW0EgO4HWngNJyCQEAxUNUTPMajOcftjPIAT0MhMkrNqkUJTcTIBYiIkU5Oc9/b2ppOJmYXAiLi/fzCbzRbzOaj0FDEjog0moW7lUQbjrAkOnMtoxsp7xKUlR//JyHBj9NGI9R7LomELNbKup/7MwJHu+5l+vq3EtsNo4OPt46pP3n6qvq7XtGZFYOtlV6arT3S5nRZcWXjA9bcnFN7s4U8DzzRPp6zqmev8Aq1/fOYDcaw2GU46i47FyVOH66/L+tPataWnpfv8roWILQ5Ay4UtQCvvzQBLzIavErqHv6ovDWqM4dy5ly5dfuPtt7926dKls2fPLhbzh48efvjhjTu3735075PZ0azLQiEgEYLnxS2OzMtuGJiaYcnD1wubkZBwmYzWbwfKxIhFcowATkD387okmQlJtL+2ExHhYKQEUIwwtI8iWe7Yvy8HqbeyMBF1ww13qjYETzq4NNxYeeGmzwmJERiQkRmIEDyDrl8gEI3Kp+QqaUJAE1ABFSeRmYAImTDFGAIRYIqcQkwxROZI5AZTULL0qooAOEkvBgognrEwEAXCEBNQ3J/lA5NMfNjmf+udWx+emR7sz37rlKdhRUVFRUXFi4hKQFdUVFRUfNnxO7/+i4RMRsTQxLA3me6kZv7kIaEGwsDEBACmWdUAkZEDcUAiWPWC6O2PyY0psuax8YP7JptBFvUneTV3z1wGO5uZqHZZjEgBxbBV259379998P0PPvnjH9/76OH+46OFAQiieRalEsqsfU+wl5khIgYOqWlSk8BZZjUnI2TgWnuJXnk7IuyICQlFFMwYKYuYKq78dEAPcnZCmkOgIWnhII7uCRBidrcPLKkayU0/mEjV1NQAXFXmJiFmFjmoartomybFGBFxMpmklA4PD4+OjmazmXSt5Kxins/KnI9GHHlJFw8Rw5E4ceW3D/YiudGBXJKhtvp2bYo27DjWYMdsfz4s1ZTPvq+tvVmVc592+wmVHqcM3Si+SYOvFDi9FvV02DL9zzeDp8Pa6D6X2mxjdp+OLwoB/VwH4hnUypsnGZxico4/Q5xutuHFcLqOT/jRq95E39ATySL0hHO/Hmb9IqA5E+pXLBVzslNNp9Pm7Nm98+dfvvj6a1euXHnllfOT6eRg/+DOnbs3bty6c+vuo08fHy1aQiRmCnFEhhf+eG3Avd7XffmLXz8hFSclUFU1AHY5c3/FG6z0AYrDkleMI2Mo7Gn13hujT1qAZdGyt2sa3PXR2fe+SjFRWy5zGmg/Y8sDZ/2eBmAMGAAbpADIUJxECMCdpAgQ3DQDvaSLlJHdXgMBwZiQGZlclA2ROTAxYoohBo7EbsQRuKfjXaMtBr4EzIAMzDBJMfmOIVBIjw+PPl3IDGw2l3mevnL0+Ot3PvnO0868ioqKioqKFxuVgK6oqKioqIDf+/X/lMgCWwtASpi7+eFhw7gTaG93kgIx+nM5mhEQi1q76JqmCSEAQNd1XdsRhZRSM5lIzlkkS44pphRjjG3bLRaLGBMRI5KqAhgzm4mqAhExM1HnYdMmWU0NCWi+aOc5pzPnr98/+KN3P/x/v/ej928/6AxagAwIGP0ZHq2PUx5kdQ6z1DTT6TTGyMxE7CJiKRHRsMLMroKYickzJHpGQVNjZqZQDD1N1WRoOITgds8OUUFAIhIR545zzrnP6xiYQwguhY4xAsBsPnfy3sxcrJ1SMrV2sSiEfs4hhJSSqna5axftbDabLxZd2xWfUGfhl4mqnN9HxNGEwJqKcbSKMJ6Jdf3y06TQy5dfFO7vGXDMKXICAf1ZsSb1Hq9nLLeu7XK8MPqYup+K5/uR/DkS3Fu16uOPXgw823ThBgG9dS42T1rb8vdUAvllg6uWGr0Pzxbt81pXrQilaUmn4vICgqbQ66Rdd+yOTqYCBF/5yutXv3n16tWvv/HGV86de+nJ/uO7d++++847779/8+6deyaAHEJKpXs9oezkMiFm0bGhf99JT2a4ZJ8RUUSyZPXEBT660Y4rlkcDh2xqIhQjMQOA5qxZiMLoi+uzrOYmzlCo5jIp7ohdaHcnqXXp+GwGRmArdtVeJ4InUjQGjIWABiqrqy5/NhqsrdHfGpkBGDPGJjSpSTGFQE0KyUXPZp5rmEwjcyCkEsWUVSQxEwGgmSgBhhCJiQPHaUwppSbu7kwiBzCTVg5mhw9n3YHp7Kh7eXrx0Wz/oNV/8eOaeLCioqKi4suOSkBXVFRUVFQAAPz+d35ZgQjSXObdorMu7zXNhJF1waDU2yeLmgGqgqq5EyQAqLnnsYUQJ5OJiOScO8mpSSmm/tle/FGfiEUUwEJk1SI3Q4TijKzSSUYKgNRlWbRd20mY7u5nvLe/+OGNe9c+vPfejU+edDI3NGBDMhi5PK9TgUbMzBxCTCk1TRNTJCYd6ISegC6C7hGIEYlEBAwIUXI2sMChPPuX1gwQDcxUPfRbVIjY47Jd7CwiQ7x2UbupmhmHUATKTir0Ps1mRojsijMzN+hwi21nVUTVqe0QArhr9sHh7PBIu84QEaknMqSwgcUHdCzdHr/qBePrTgc2ZNoaBY0vPx0NaIynM4PrgsxNIvfzxmeu9TTKXtzy6Wlo0lHnTuJuzY/HaGmlDxsYWh8LsNd0nxvuvCfh+cndNeJ8ewdO0+7oZNs2rz8FHMPirny0yYD/9J4j8Lh3uPHpiQS0DWW3rUnYCe/6C8Za26NVqvU5wI0XaxtwfQ4RwAxVkQnAVLIH0ADi3t7uuXPnLl587cqbl7/61TeblLque/To4c2bN+7cufPwwadHs0XbiioYICJKzuo+SH3nig6ZeCtLrsOyjgEiElN/M/L6wLKYFSMjQAS1wdMZ1ua0N++A4uU0UMalPLGvIfYy6BI7gr1ieqm8XmqffQhL+fPKugEBMEAEiIAJKCFzL732zgUi7i0zEA2dd2YmQrdv9lkeZokIGDEgNhwaptjbRFluES0wssdCMTFTDKFJDTEhk9umqFknQLHJWeaL2dygFVsIfPxYL0zjhZ2z//C7310/JSoqKioqKr58qAR0RUVFRUVFwe9/51ePTA6Rp7MnphaB9iYpIkI7h9whmKiK5KzOoI5DrcEzDRJxTNHUXE3GITDzIJRzo0wEcvKMuA9KLmpiYw6iulgsOCUkbrvcdlnEMAQLSbn5+Mns+keffv9HH916dPDgaN4piZEAQU+0GMCQt6qHGUBgTqmZTCbNpAkxFl9NWBLQthnYjgCIKoqIkUhEDICIVEpGKSLkQNZrlnH5ohheD4SyM/LFRrNPe9jL1VBFwIyI3ayjSKRDKLyEaQnPFnGNmqoyU0xpd2c3BM45Hx0ezWczabsskp1GUekdokccyhZgz/CNQ8zLvOGS+7CVv32Bfn5P4KC3SIPXm4F1VudpeEbF6LKdEQ/1OZCssKxwU7G8WXZrJStzPghK12ruvz4DBW3LSRtXMO7FWssbU/aUGd/wLdhy0LZhe4WnPGAbbOhoNo9t8BmI9aeVOp4+37I08DkKvTdxLPsMJ0mbj9npJAJ6de8tBPRmT1YJ6C3s89rrjVY3F6BMiV1um0OMzWSye3bv4msX33jjK5cuXTp/4fze3u79T+7fvXP35o0bt27dvH//gSgwJw6pOFWYSdeZKviCjEFhcgGIGYjW20fUkcy5WCQNSWbL0p8UL3/CZVgJjmam/5+vH/omRNTl/adYcDDT8mY35BsoYzfnnT2VX3/NL+c8rnwHlnD2uQGMQAkpUfA+opU7W+gpZkQDNARlpsDBbzJl4J4bUQ0BAmNgSsxnJpNJCAEQyRDFtIsBU2RmCkwciAiZqYnJV16zSCea1VqMiwzzeScBFXVh+Aqdfzg/uH+4+IMPPlg/ByoqKioqKr6UqAR0RUVFRUXFEv/kO78augVpF6xli5H55ckkcND5jBFUJee86LouZ+dDR/6YKFqMlpkZALNkEVFVACAskipVE/GkhSCS/ckfELPknPNkZ6pmhwcHHBMyi5h69LIZECHx3PhJS/eP7M/f++DdD+48WcBCMQMqkAGZZwMciNFCoZZneuYQQ7OzM01Ng0zWkwjOQbddJ6rjqVBT73wgTiEM7p2LtuvaDAAxxmaS1GwglKEYiBoAcMnEaESkql3XETExFb5CTUUAkZicVAYDDuwmHiUvoioCMlEMwQXRPv8us0PEvd3dELjrukkzaVISkf39gydPnnRdq5IBrI/jHhxXN0n2tUSO/cFc2QIblOYGP7kSz38spfW54FlNkhFxCJkHBEQaguuP2eH4urZTfTjW0/cyxKfuNpyfhVxeMv5jxnAsY8XBEgDNtO/sYCM7mAyU02OlrdXxrohbVz/bYjgA67X1baxOQ7+kc7J0eVXbPB7u+lk1HDjnAzfrWu3VqU61US1bKXgbDWSrYnhtUKO3J5+Xp/wi4LFvtnRnS4MjqhSOGWLZtP3obMB6TS0AbuPcEUcbN1vSjS2w3m7pi4EpiJ4999Jrr1/8xtWrb7755usXL6aUnuzv3717569+8M7NGzf3Hz/OnYgauOmx20sMY3Eyd9QxN6Bea94t+HUghNUQgZi99wIGKqYKSDAYeXgGVPfKWPH5WH5Z0KC38tA+5KUciMBEhFaS+Rr2zLIvTIp0JgKmgOSjGM2Tu20sx4AACBbdeQMoACbiJsZitg2GxWxbwfp8ve6yDWpmWIhycBtoBEghNqlpUkyBE9Nu0yQiUCU2YggMkSkGTk0kRgNtF/OcOwDIXe66tu3ajIRxmjl1ispNh2bzedNMAjc7OK3a54qKioqKigGVgK6oqKioqFjHP/+1/wCRkTkqNiGcm0zP7L4UGUxFRbLkTnLOuTy/q4qKW3Coqog6IaCmkkUka88Jm0c4D8JZFWImok6yiKppM5kY2Hy+CDEiBzUEIjdc9sfxhcBCaWbp5r3H79+9/97NT+48Onx4lAVQAaUwGZso9BwRxxBjSs1kCkhaArFLyihVy5IHZsHUVBUQGCnwkO0QVFXFtXVEzB5UPZDXZuaWooPWzdM3uZUHIBCR0xYi4r0SVesJaOrFelaUcQaAKcYQAxHlnHOXeyE1TpqGCLuuizGlGImo6/J8MV/M5/P5bD6fgci6N/DarCB6wDj2swTouaW2iJqXQf1PUaVuIaI/ZzzTz7f1bnxWCfQ6lo7LW7s1EHiFjsIVIelWChX7IP31lgCstw3oz/RNb+hNIe94dWDlo0JArzW/2WrfyrG0fd/UVpJyiWc6M54quv5sP+KHy9Cz7XZKKfhK0X7to393zDRsKo5Xyp043LXT6bhRDcVOO+o1tn2jPysE9LbdNylrABiWBk0NDQmblM6ePfPqK6+8cemNi6+/fuHChRijZLn/4MHdux/dvn374YNHR4dHkv2CjQqIyO6bNJx7YKZmrkMeLU/Y1umw8Wh6P2jwVTs1MB3Uzn699Qs7espc11YTISJ7dlm1Qb88CJex59+pfPVNVcWXMVVNireSlqyD49nFUTeXNhwIEJAScQQMSGxAZgQYmAcSvxiP2HJHBGP0zhgjMFEMHBAZMRBOmmbSNJEwhdDEGJkYAVSQEcjA74KmZpZF2ixgHYIyIXtED2GY7sxbOQDsKHRGBAwqkLvf/uHt40+MioqKioqKLyPCX3cHKioqKioq/sbhl37z//rd3/gFUhNQUZp17Q7Yzu45kFalmxCYWdZB8ytdlyVnMyx8tIgO5LSqC4RFREXMAJHdMRrR/Bl+3rZqioAhRQPglDgE4mCASIxU3JBNZZJzVlBqzp35ysVXzjWRw80Hcm//cNEuRGSd7RiLMd3FIovkTjIgI7EaaG+A7GHHrh5DQADCXn2GgKa9wswJ5VAqVDMiNrTe99MAIQRmoi5n5+s82aCZqYiZoQvwiidoIZrNdeJE2NPTvTrP3aKZmZGIzNgscCBC9y11tiLnrKYxRA68F/dSShzYwLTrVER08BW1JW3kkkOjPgXWeLpOxprEdZNCXTJC6xV+dh3oenWnICG3c3qbW0/RuZU8ZqNd1mi4TVtrP6fURnTX1o6WCbTtIxuoYBwfyvXDtrnjyZM0kkNvZ5iXFB9uGdp4Vrby4KsfDk2d2KdSHrecXSs9O2b7abDs/PG8+sY+y+6Mmt66N668HqcBXTp0P+XIodOhTz/H10/LcizLaTkIotdc4E+7CjAcVCzfaBvePq1nGwVcS9x/W9AAOYVmks6de+nSpTe+8Y1vXLr0xtmzZxdt98kn9+/cvn39+gd373z04MHD1ExjSGkyKU5HWZGYiVdr71caPSSndL5cZodSqmquqy8eSOV6u9bVlVIjAtrDevzyTESEpAiIAgqiamaEAUcnF4Cb/isYqEmht3PObbfS9XJ9GM88DAfJDyQBJsQdCozIgGBgKmbWiZSRmoIpASICgWuckRHNg5DAYqAmhmmTAlIkDITTJjUxgubImBjBBE09R6MqtF3XdV3Ouc1d28milSZhE7mJgZvQTJrUpE4NIpqyqqWHOe8ZpPDbP/zgKedGRUVFRUXFlw+fTTxRUVFRUVHx4uL/+Af/cVDmjiUJ/P/svUmMLUua5/UNZu7nRNy447vvvvtevhwqs6oW7GghJFpIBUXDqtVrFkgsUEksUDeiG6Re1Rax6V4g1Bs2zS7VoKaFQE23OiVUIBbVi4IasnJ6w53nmM457mbf97H4zP34GWK4970EobT/y4wbccIHc3M7HhE/+9v/w9CGuYGk5clh28xnXtCviTEwBygMNzKxW3p9cXETIzNnkZxzzg6pAYAcBJup//GfVMxTlQOJ2arviRiQRFQ8gkMVVNGUCM0gZVVqVxBenuefPXr5p7948he/evLi+HxhIAB6BVpBRCaKyJE4cBNCCDEEJ88el1HWcRuAmeNjRBxtbjZs4CjZqzCJqC/XZmYiBDCHETBkceTBjKxmRMTMTGQAJbvDTFWdKTOziuaccbA6T3JDEQBAC80qhaJExgsjQiJP3mYiXC6Xi/Pzs9NTzRlUAQyQgAgNwNRMANgZ+xqI4k4cdol3gJFGrXnaBO9vd/OWa3NEtXCtX772sMZtZjv1C1+m/Wfbs891APRkvT+gjQkDGxbjtb10YHX7Qh0Ge+b+hozuza3vr0fBpqF286WNPWxr58uvcA+r3I9nRxi+7o0N17aNI2DTg78LzHcP/L6u5G/uZ78mg94Ti3y9nfcEN19ZfPNaf6N8kz9kvqGn/EPaTCUwxr260Mya+w8++uzzT7/7+Xcefvrwwccfr7ru3bvjr7969MWXXz1+/GRxvshJDBCRgYiQDRAMVBR2gmEQEYl8focmTSmV/yam94FTlzvqCfuboxc8UZqIfBZQVb1Orek6xRlLHs5w/JJ3xENnWHkWmGKxVquZWMnD2On/NYDG4UlpBEAABMYADNggt0Q82r3L2x8QSkFcv+zIHIjZ6+EiuAOaTJrA87Y5mM3awJE5MBAYqqokzVlSNhUE4EBIpGZd6gEgMLWzNjQNhzBr2/msnTcNEinA2eLsuO+XSAtRWp1ZjrigHz96dMU4qKqqqqqq+o1UBdBVVVVVVVUX6l/8Z389YeqktxAlAampdg3khiDGpmliCJEDewGkGBv/0xhK5K41bdvEOPxt7rZOJOIhG7o4oLMWTxkxi8qy771onoipoRqYx16IEIKK9F0vyBnCudDz4+XXL45/+sWzXz1/8+Tt6UKsU5DLlo6j/0WPxBgCxxiiA2j09dRZREWc7aKVddYlTLR4qMVGAF0iOEBNCb1AE5fCUkPyCCEBgA60PeeMAF5m0AAkSynAJVJSQohUTSQXr7QzcXdPIyKSc44hjGGdbkzo/yExxxCaJpiaSE596lervlv1XadmAFRMkaYFbgCsGfQAZSZdNgRMDOhwA0DjxqaXaYdsXrXt9BbiGnhufB8v2GGy6+4XOxz4YiPrzsE23KabyGoPWd3C8FuvbyLbrRPtbg0D6TZz0AYj87q0Xye7X8NOu3OoyRDY2GTPZhMaXnrEYGOUbBHDnRaub8d7Q+hvyqCvPsBVXXzR3dw7MbB13I1M7e1Rc9H4+YZ/xdjm++Eb0+edl3c3QlBARYAbRzfu3Ln98cf3P3n4yScPH9y+fTME7rr+8ZPHTx4/e/70xavXb49PTlQEiUNsVYfZnP3588PxyZ8TOJn1AViPpsmoQhwfeqY6TuOtj+pPWyJfoWLmBQ5LHHuJJvdZwIFoQ8HcZTUMmoEzaA9fLktapJiV1+0eHj+TxsGQjsTD/wJAQAqIvlTHndTgSdUAhP5TrRQejMyBmYlDoMBECIzGaE0IMXATgsNxNJWcNGciMxEVYQCP1wgxhMBEGGNoY5zN2xAYEJiYiIkIm9miW705X3Sgqx4XKw5hxbb48Z+93D82qqqqqqqqfuNVAXRVVVVVVdVl+if/6b9tQKaWQVNWlD6AyvJccw7MgzvYzIw5goGaOcmNg0IRMwfmEDiUyoSM7i/OOYuqgRGxmqy63hAMUM3ziIvPN6ckkiSl1K1yli7rIlmmpsfmyevznz168X/98qtXCznurRtrtI1esvUf+FgYNCIwIgd3IyMHIgJAL67IzDQpXofoOZuYc/b8ECgZoCQqfsmOMwhRVSXLcE4EACQk5rJ4vE/eOo4RACQLEiKA5gxYIjhsMEQjIXv9Q1UVgeEcAGCDXW5kLiEELOBeECEwHc4PDubz+Xy+XCxOT05OT05Sn9zQV1boT0HygGN24yF0k/kgok3KYu1B0PucuBvfmbDaqTd6co7dI+zTTibCnnOOsHdv7MXQARMGfTHmXqPXsZOm38Kpz/Lik43UeHeDrbaXk003Le7RMaplMNpfR9fZcn331w7mPXutAd/OwXePsOdduLHnuFn58mIuv3efD0XPEwD7zf8emN76C7Q5FbI5GkcAfSXqv/7tvoa2OnDry/ETuuIAF4i2WoqGqMQQY/je97/3wx/98Ec/+uHdu3fm7WyxOH/67OlPf/aXP//5L549fZFXGSkgs4oAEYVGs5go+NoURF93spbt77jS+L3fRZiUYDVUgWF6DfzucIDhp9uwuwIoePA0opkRopeNhWHhiJkZYPk/aDFBey1dA/MIjiEGemx6uYh1Tgv6TBcjBsAIFgADYCAk8Eq7YqZYgjWIARkhDD8cCB0ic2AOkWNgJgyMkSgERgRT7fsupV5S6vskIrO502ach9gwM8GsDQfz2dGNg4O2bZvYRFbJ3WqZsvRJVilrOz/u+i7wqgfoo4Ikgf/xpz+9bEBUVVVVVVX9ZqsC6Kqqqqqqqiv0j//m7wuIoQCwCdyc87yZ59XKVyS7zVYkq3ixIhMVVRMt1ZBgYhD0MoAiWR3CMiGRaIFBIUYD6FPyP8AVnOgSAKhqzpq6FaHdOJynlPqUFThTTBBPe3t9np6fdn/+9fMvXrx7c971ajIgpi2gaI4PwL9HiISE7fwwxMZZMDjeRUTA0QG9Jo6jb85Tms2A0B3TvpS74Mk1hhsRK5Kv6Xa+TASIDhDNY5oRiSiEKCopJWYuJjtfWm6lINR4TK/3GEJw/3iB5ggAqCI59yGEJsa2aWJsiKhbLhfn54uz89VqlXMegOna4jzEp66rPrp01+yK64tab1s6dR8KHunk+M8wLvYA6D2m5fXxN3UNAD395AoT68UAerdJOALa/cfaooYA4OjKAEAFAIG2ij3usRTvct7J8crUCI7du8eCvXVE29cFdslXG+2yyzpyMiOxTaY3N78YQO/st6avuzv5FV/9i/wusJ3mzezptH0O8C0T+nhQ3Bwzk3Ptn0/ByRgenydjQy+zfe8+Tn7NmkzYlX/e+48m2r5t9vHH9z755P6nnz785OEn9z76aHYwW5wvXr169dVXXz17+uz1q9en5+d9lxCCGSrAEJrPZmYi5j5lRGT2qgA7N29czwFlohHWIdjDNsM82xDdjoRMm280ROLglfeIkJGYWTSrKgf2HwlejRCHgA+DASzLOCfklQBNRUzUHdBgCsMky7CmZBtAYwHQFpEiYgCIiBGIyZfhKIAhApU6jMiAhMiITEiISBiDV07wx5Ohs3JCUwVTRBvmOp1WU9OGwMiILXMTuGU2zYQ6b5tAwACzNhKimiJH5eb4rHub85JY0NJ5BFJQ+vGf/dn7jpCqqqqqqqrfKNUihFVVVVVVVVfob/z9f/6P/ta/CUag0LQoFA3x6Na9gACaVTXnlHNvoqaiqinnlCVlKYWc1EoZwiyImEPKOYmI4xsDUEUkDiEAduAUh9AAxICIyCtNGRpAt+oI4WA+K6kUoJYFIM2puX/UHB4eJBEkjK9O3p53Z/3Uh7xmWe5sLs5OM0M1Q029AiCz27qV0ACGclloBqqKAAUKD8WlDIwInSwXnmtGSMSkqgaGgIRoAFnEs0lDiAamogaGSBSilgjsAhxDYNJSZdDdar7kmQjVTFVGAiWqABBCyDmriNNtQCBiRTQVABDRrk9EIYTQtC0hNU27WCz6rkspSxYRsbXF2cHIGKO9E7x8EQicfNOvuryy/e/6PPsW0k9Wze+FXReg3s3Ptpjgln9432G3v7e70fDKRvT18HGHNg+W2onfeV8LcNLa7aTm4fMLegJthGoGgEPRwmm79nLb/QgRN7tx13+M01mG3VZuyTa95tv24ov23AeUrxwIZvtnAC7Whs3YcPu2I8LkkBtHviCuGyZtvGoGYLsLL8L4l1/0pTT/16HpPNGWRmQ6Qe9IpcZpySAiunHj8OjG4dHNo4cPP3748JNPP33YtI2IPn/2/Nmz548fP3n0+PHJ8UnuBRA5tMyNGYh6uAyiP7JZ1wCaGExNxSaPEkRE4kkceuHLw3oPRCgLfWCAWAAAIABJREFUdEpCxxg7hEjM05GEAERkar4VlWlKRkIixjXbVXc0+4SQ52ygCnhIEg7fEDEpFmgowfHo+29C7/XEEqHbnyEgBAP20xmAFac1ITASO4YGYkIH5YSAzqnLj7cCoJHIgCwX+txwiJGZMRAExhgdQENAaIhmkUwQDKKlYBiIGoIYA4VgoXlztjqTnDgkhLiaWUw5VfpcVVVVVVV1taoDuqqqqqqq6lr6R//J7zEjGlFDEcO9wxsHhwdkYgA59ZJSE9BMc+5T1iSSsxAxE4GBqOSc+743NWbqul5EmCklSSmLQGza2WzWdZ2ZhRAMQQ1ElJl9jTMzM4fT0xORfHAwzzl3fb9adUlUDblpldtE8TjRs5PlXz569sunb5+8Pl+Nf+4jISCaudFNTHWNGwplRgrETWxijDHEIAa5EGwwUxVFgBijAQwFBg3AAhMgqpqTaxgg9arrPKmjbVsA7PreAAixaRoAENEsmZnbph0QhoGpeSlCImb2MJDSRMQQArjPbpLk4JQ6pZRFRqs2MSMAqI2+7BImDXBwcHB4eKPvu8VicXp6ujg7Xy27UhcLRq+gUxIEYCICIluXx9rHobaY6kSjEXGy7WDWXa9q32euvFZW9DXp2xaL3aXqpWFXHAAcZU0PODDkHb8rjqZ49TQVmiQjg9OkKaSdAuirMxY+zAS72869Utk+PlExll7ehgtuGW7su3l1F8YmXFvmUeaXaM/tniT0bFFd29pu45sbBx0vamP0Xnzvhjcy7TbGvJVg4+577cYXpwp9sPaD7p35h4tPMnh2CcxAFQCRiGMwFZOsqoDWtPG3fvD93/7tH/3u7/7OjRsH8/ksxvj8+csvvvzqT//iz589e3FyfJrVOMT57MBpMFEwACsBM0PX7UwIGIDBergiUQxh49vDZ6rGTIgoqj4p6GR543jryylXPUQfiXrkMiIOaHd4YCqYeDS0mSIYDo0e5zfNHFJvjlKEyQPBhk4s9QwRoCGecWQzNiMtMSJUjMwEJgjASEzESIQUiJiRyOOZTFIPIkzoP0CZqAmxDQENmKmJ1ESOTAENLAHkGCh4rULRgBaZ2kgxIIHO2+ZgfjA7OGzmB6GdPXn99su3Z28yLCWnsOQ0j/38H/7Jn1w4RKqqqqqqqqoGVQBdVVVVVVV1Xf3jv/n7FIxIKcwitXePbty5eRsR0TKDomUzNZMsmkRFTbKYCCK5BzqlbGbEJOLJySpiXtIvxKZp2lXXeQFAw/KHvCdgpJQIKcTQ9z0ANDGKSt+nxXLZpySqgCyAncFJwne9vj7vv351+vXz40evTs66lAFgnZgAgLCTm4sDNQwxxBAjx8ghILGK6UCICJEZCy0eLGYhMADknImJaQwVBRlAHhEDYPYqhcxMJKI5ZwBDJGYuMR5ExdNn5tBAh3hf/zgAaNjyfFJJplbnzv4tAmQiJ+CI6J8E4ibGpmmIGQDMNHWp77rF4ny1WvVdr2WFuA22Qy5YGvehrm2uN+ViQ0PBpmHJiOOBNq3Eu4TrChY5OqsvcYyOR8Ky+B18IoK2LMfrxm5p37GnMG631cXAiGMGy+TUsLHGfxfqTbJqtr538TV+ALG9hrbatkHldr3QW/d8m+Fe8bv2tFMGi2g507Xauh2vsO8Mu23YSizZ6xaf4t0dV/2G69lw/cJF7bnmjbp4LmefA3rPiTybGABoePtfpmsC6AunnSadgIAAVsL9WTUH5qObR/c+uvvgwceff/7Zw08e3P/o/mJ5fnJy/Pz5y8dPnjx9+uz1m+O+zwYoBoDEHFQMDIcHlJVSrjZ6mv1O+BPZb4utWzNJSrLpQDJTM0ICLNH5iOPWWDa2SQKzlfiX4SnvdmY/Iap66IafWUtwhhmClYBmFTMP3CjvCB3M4Bs9vwOg0QDNECACNsQtRwYgA7LCxhHUrdheJ9B/2JSlOmZehoB91tfcIo0cODAxckAKSJEoEDIZoxEIWg6okfFg3jRMgbAJsYmhbeO8jW0TiICJkdiIM8a3Z6cvlqvT3pYpH58yzjprux//H48uG2NVVVVVVVVVg2oER1VVVVVV1XX1N/7+P/+f/s7vEQYWyZjPumWzag7mN2bNPEDWDIgQApWSggCp7yVnpEIT3NKLhCrqcdEqpgqqyBxCiLOuF8lm4DWmvBAfAPZ9ZwDMHGPwxdQRIMaGQuj7PqXezHpRy/kgEoZwcNAezJqb87ZlenG8OO76VZIkBojjeulNWeFqmlVA0AyMkJgjkKF5JCc5VOSyiF9VTU0RyeGCqSkoDC42GAiDiBgAACEDGqioiKgKIgFoSupGZoDBLjtobFvJfS4g1UmDt8G8XZKzWYE0qmqqBGAcZAKgzUyZs+Su74Lz/rZtbjTz+SzGwCESLXJOkrNoRq/9iAju3TMDvAAl7gGF6Ah75JEbhmFEnHIrv473MXKuzaeDjXivo3kUIYKZJ75gyeAGA12bTadHmNqEbTs9AgcAVr4cLZYjIyvZrtOr22zexU1dg9KNbca+mYLayU7X0nt27/ZVj2+ZYY5hB0kPzvC9760LmzmG8A5bbpqjr8Wg95qFt06/u9N6CG0caXtHvfi7V3/jvTbZ0SW37LK7OQBoHE78zSzSl5y0vMFxsA47njVCbCK37ezo6OjBw08+//w7n3326c2jGyGEs8X50ydPHj9+9MUXX714+er45BSMQmxjM0MzVUg+MalIQZ0zqyoMb64BQlt54yHue08MD50t9/r6MbQG0zgWM7TNgTsmtECZjANCRDS/QofiJbHbHEDjeEoDz1l+32UKaABm5PQZqAFqAMkd86iFmXu4kSeQlEgRKCEkCGZGQ04HBWImRgzMzBSIWQ1NGZHRGIxBCYRAGsJ55KM2tjEwU9u0bds2bdM2IQRSAwFUDMuUXxy/ebPsVoR95sev5WgGtmp//C9/8V6XWVVVVVVV9Zus6oCuqqqqqqp6P/3T//yvASGRCLVgzc12ftjMKK/ActOEg4OZgZeJCv6HMcfgBY9GtNr3PZg1bZOzpj5LNkJmCklyFlFRYgKAlJIjQwATkZRS1/Up9UmyJ3IgYdf1q+VSwbJKlxLPD5WbRS+94jLBq5PuV8/e/uzxi0cvT0+XvTElVVXb/fGPRAhgCkAEREQhNLMYW2QCRDQUESuFE5mJ1CznnFKiQGoqOVO5xingXjNO0zUxcXtsqSuo6nSbmBEMTHPfmYFTeyIiJhUxAw5sqqo2uufMitnWcjZVDKHwERU0A78FiKLKxMQEZswcOHR9T4gH8/nh4eF8Po8xdF23XCyXq+Xi/Hxxfg4D4S6G6L34achP9e4br/Qila1pTND+cA3Qc33CSxh04aOD6ZVK1+34rsuFDFR0OAPAcHXF6riHjdpoAfUvEWA6DHZSF8ZW7b0uP9fAwIop2NaAa7rn1b/H7kXCl6R8UKletpbqGCCwJ85i7SEdjryNlctmayI3BlhvbWmmm51yxdXtPdG2Rh/qxnERrqbbun2H9sVjbxPwacdOruzq++T9c40NYTTUrx8vW61C2HZAX9Crl51t7Ua/KIKDiH1uDEEBFNDMdD6f3bt77/Pvfv75559/9vl37ty+M5vN3rx5/fTp0y+/+urLL7989eJV13WqZkBg7InbvsgCCu8lRJ/KGaqz+oRWeYQU3rpxFThp85Q+m02miQymN7A8hAcAvadPqExvMZeCfSWCQ8dwjdIQU/S5CjNUNVmngpS5yX3zAKNXu7ibDQisAWqQGqAGMexMBQEMmR7l4YeBKRAVp3MgHpbRBHanMzJzIA6ErEI5B4CGqW3CvAnzlmeRW8ZZ5BsH8yYGJFQDJI5N0+e06vqzxUq4XWRZ5twTKnDC/pfx4a2zd/27s//55z/fPzKqqqqqqqqq9qkC6KqqqqqqqvfWP/u7vy/ABqhKqhSN26YByRHkxkErOQMY+VrgSCFGDkzMYKampiY5A0CMUdUkqwogElMwL+okAohmlnJ2bCBewjDnPqWcs5iSr0EmyiIpZ0B0by+3MyPuxdQoKZ12+ux49fXLs58/evn49fGbs65XzfvomxemskIsEImIInGkEIhDYMZSZrAgInWncSkgqGbg2+Rc8pQ9chQARNSgHBEQVcRL/o0Uw0sMgr9koqJESBTUFBHHMGgnSgOALpsXKuJO5yEAhEpSabHPWam7VbAUEaWUiXDWtjE2IbAv3PY2pL5fLZddn/q+77vOCnbfWcu/tgyPGBr3JAVv7VRskjt0cvywYZjetxVMTcrrVfP7fp8bjqPD5ePgT8Rt/riJn3DNszYPj8XiuNGGPS0sGKiEfiDRXt57gft281IGVrtp0Hw/fr+z/cUAeiioubG1jgEmgJf+5lwaerkjfQpycdrXI6ybjJD9zcRhk2v9Gj/y7sJqx703d9/D+sZhv54N2G3J7v3ac0ScHGW/0FMcLttkzykmr26fdYr81xtstva6ABrXL052HiLmFcACUxPp7r27Dz7++NNPH3784MGdu/dm89liuXr75s2jx4+fP3v28sXL45PT5apHAOJAxGY0hHijhyX7QCPGwWWsZQZhbMI6xWesIegVaodOnsxzIABSKRFrIr6upYwyLEeYvrsmdHqchQIkxokAPFOjPMUJwOf8VNVUQBVU1yP5AvoM68kcAzA0YICGKCJFoGgQDAgvJNdDhDUyAhEQIDMyIRMgGIJF5sDEBMwhEAXCYBbN2hBmMcza2MYwb8PBLBIoqcaABppFc/bCjrhMKRtlajLgImcNlEFjhBW2S4xv+egnP/nJJaOnqqqqqqqqalcVQFdVVVVVVX2I/pe/+++BGpuedqGXbBkYbBZ4BpJSr5LBIDYcmhCaEEJ00An+97MBIpQQS0MDHKxahB6yCaZmWbIZmGnXdSIKYKmEeBCAOFd1/xgRiciq6wDREA1QDZPgMtt55pOefv718188efXLJ29Ou36ZRWzf3/YDYtayhp0AGDmGGJumaZqGQyBEkVyyRBCRsE+9urM4BERMKauVcoVMZAApJQPg0HhxwpSSqIiqibqFOcbo7TcVMEWkwBxCyDkbABPJRiLHGBdSRAMW8X+QiImwLBW3kVyb6bQcHBGFELzEVt/1B/P50Y0b84M5IkrOy+XqfLE4PzvPqZec1KGETeDgdoa20+edX6t2USROPttAylSYV7E67t6fXbo9Nbdu4eDJQUQJiWIAAFPVlIHIDebrA22aIDde3n1ttxUbF4hIDGCmAuCh0zymsmxsuP5kwKFTejnt5s1k5PdKfl6bQScxBZcg7F1b8QTg7jvuVovfV7ZzzUMb1nXbDDZh7uZI2HUAw2T74hgvjtHJmNmZhVj7aA0ADMcI3zXBn7yBRkS+21d7tDM1Y5OzGZTEmm8CoD9IV9yx4vCddLhNBw8R+txVjHwwn908OvytH/7Wd7/7+cNPPontTNTenRx/8cWXv/jFL588eXJ6cppTwtAyRwqeD0FaXOaEAGqQRVUEzDjQZgDztLXrCI6xoqPh4NAfWjn2EgWfXCPJHq9Pfg04WJp1pM8TagxrhzKMj9fxSeuPUzNAMEbQrCJZJHlBAzNDWz+P9j1BhgOCz3YaATDijDggMSCLko3hGuNeAABMxBwYiclnihTBEJTAEIypkOgmhhh4iODgQNggtUjztpk1sYkhMMXI8zZK7lPfifQp9X2XetGUtc+SiZXazBGaiEw96/Kd3TqigwP8b//op5ePm6qqqqqqqqq9qgC6qqqqqqrqA/W//hf/zrtVerM8O2qOJGPuRXIC6YMZiEjqOVAIzIFDiDEGJuYQQgiMSOhYAJEohhhC9MgO9/x6EK2YjuzAM6OdyYYQRLNoFhHnSH3nFJiyiIiqgailpMteknHGeNrpi9PVo9cnf/aLr754+uokWTaQzcvZcbQSgEdtEhFxiG07u3HzBpakW8cv0Kde1RAxhEBEvkRarZRPdCs3EnFozExNVXSoEoZmJqJt2zBzFjHJprr22bkl0BQATC1LjiE2bQNIZqqqZWH4WmUHIjI1kewuOUR0CzkzmYGqxhgBIOfsu6kqMwdm8sDQEA5mc0Rcdd3i/Pzs/Ozs7CynzkQAqYA7X2ZODO4EJALA7aX6CHaJJxrHRJI1krnUAb2564gW1y+Mr0z6xMqqfDeDg7lhsxgI11vtB9A75935xXELWo3tm7ZtB5EOaHnPCQuLnB4KzECHoPBicn9fB/R4WoRNmLenAesdNto7uRaY2mP3HeEyX/pF54QyIiY3xYN0bZiWoIvG0p5gkOEIhmADI95GgluwGAE2bts4xK4QbjLo7e61IZZ30lzYvEz/vu4bX3tPeL3NrqXRTTy+hYYsDBwbSlwiaAB8LKqoipkAwGzeHh0dfeezTz//zqefffbZ0dHRbDZDpJevXj15+uyrr7568fLV8buTlFVKeAQBEceAiGAg2fEzEgUcigQiGPGWmxl4/axTv3oxk3GKYr1EwxPzDXHwUI/p1DZOQkwYMAyAe3+Prm32Vu6kr+KRkg1ihiKjU9vAX7z4WONcCCIhECADBqKIFBBBFb3xQ1oIIfGwjAWGSVFCZEQiYEJGCwiBkAmYIYYYAsdAkTkyx8iEGJBiCJGYAa3UQDAkMtCUUpYkmkXFf86pqohlgeboVidmMQpCj7q8+535yWs4WdbYjaqqqqqqqg9WLUJYVVVVVVX1gfpr/+U/+wd/8FcablISFs5UeDDFRrRLqtQL5QyGiCskwiF7lYiYiJk8+zgwcwhMbGCEyMwhRGJSU+YQAjvhJWYzRSI1MFMxKGkK5KXlgCgEIAQVNTBFJmqCAirx4Wx2dDi/c/NoFvjm4eGvXrx9fbY8W/UwVI+6wKqmYGhm4tUSQXkBIUZmJgIDT3wuXr2U0nShttfPKnTVwCADbBhhvaqhlYRfMx3AxADa3I/t1wgERMi+bt35CSINUIY8wBpMRJ01m6qKuufacYwf1ulRcPO4M03vWIAkAiLMpGY+YRCb5pAots3sYN6vVn236vqUcjIZ0b0hEtCYULzlBgWA7Tp+G707IC/AMVd5Ygvev8/Wt6am1b07Dox77Y2eOE83jLJX2WgB3LC4eZgLWznsPn7cbPyQkLABT21vB6DBEF1SKOF78cftooiXCjc/XIRgN93rGx01+lSvrTVR37l3TgivgOa7odyTb+1J20Dc7Omtc6+H1HU6bM914tYGW5nn/kDY5OHfnqn5g3WBdRtGRFvq7qmZMmPbHty6dfPeR/c+fnD/04cP79//6PbtO6dnp89evnzz5u3zZ8+fv3jx6tXrrkuqhswByQDFzICQAwCAGZD6UhgaHL0+h7bG4kO7bE3dEdZpJWMn4rTJZkBEDosHR/96lgIBef1Wsr1jyyYP6/UGE0t8+SgiOY3rFACmt3a7HyfvfKDhfwEwAgZAtnW+c5neKc9Fo5IjUlrOhEwYyAOgIRAEQkJjgsD+HxEYmoCCqiUzkyCAqOCzswpAjKK6WC2zioIil5+jJmKAgmGWBSgkST3imcCN5cny5r2f/MufXD6Iqqqqqqqqqi7Rt+UgqKqqqqqq+s3Vf/cf/d5KcsoaGEMAE8MsmnqVpKqSc0q5KPWpW7kBmomIeL3CeRAhtm0bYlTVEAIHVrUQ43w+d39ujBE9lJk8aZqZ2QxUjIgMLKUMBghEFAxBTJNSxig8O0326PXJ//l//8Vffv388atjRVMDMdA9hlSc/A8K5kBs57PZfM7MAO5MNVUTUXWbKmEMMYbgVjMtmyB4OyeFCkMIAKAqROQogxAIgZlHsuwQxLtl9C9nLY11B7l7xp0vZ5GUUkpJRQk83ANV1Rere1625Ny2LYfgl7T1qxACMhEABObZfD6fzdq2YaauW52enr5+83ZxeppXC0AyQDCjEJBYU3JX+HYX7qu/N5xp6NiJ7/UiK+tFup5tec8xd2ORr2t3hTJYL2vVpRcxiX61jVc2tin/jvMTF215pfaGQuzJA9nTBpxuabu4/NImbe14HV3Rqx8aPbFbQ492r2LYZnIWgxLscOmpJ2T0wk3WvuLJGTe79/9jB/R47OlkwvDmJSvp/cMDw2YHs4/uf/Q7v/OjH/zg+5999ul8PlezxXL105/+9Gc/+/mvfvXF+el5Tjm0zXx+OGvnKYuoKaD4fBOyAZiaiRBRYEag4k1WEVPJed2s6S0pbNq0zMgMT2YsgxMR1esbEvrTMnDATe88EzHxeGCP4NgaEmaWRaZnpnFxQHERG6hqyrlf7fTk9mNw7FW/RvK4IrTg6BmBfakIqk9nKpkPrGDEgAEoEDETA4VAMXBgikwhsHufCQ1NwZSGSUnNPagQYe57yUKEoGBZPRGIOHAgA+v6VTI1wqZt1KBLWXOmEHvD+c2b3LSrDv63L7/8rft3fvny7VVjqaqqqqqqquoKVQBdVVVVVVX1Lei/+Q/+jXRwHLujNjSHkW7fOLx5dANMTXJKOaW+7/uUUupT33dZslcU9GwNwmCApuAZ0Gbq8dAi6n9QZxVADByGdArwrGdE8kKAsWmYGLRkTagKUwghhBjVIImoIXLkZt4pnvTp+en5o9fHj169+/rZu+Nl3ymIr+LGvUCmYI7y13sITpIdKQ9+ZBLJHtbMFJh59NAVOxt57ggOi7iNvSqjikczqyqh+WGnYaMpZafPMQYRzSIj1bV1uAQgIDKZqmRREQBgZlOBwoW9CSyqOefBGb3Hx4sIhGRmHMJs1jrfn7XRdxERSVlyf3Z6vlgsUt9PW7L7a9UuUrTxlTWAhsHrun+XS7QNoNfjY9zCpv7nLeq3mcJxLb55LZyN21vtEkwvjTYedDR97m5ZjOo7n19T/z8C0HuP6Vb9Dz7UnoMD0GVm6jVzRNgG0PtOfx0cvDdvZct6a+VQV17junM2bL8Xtm9E3PtG7p5JqPFiEQAMsRh+EWA2a2/fufPwk08+++yzB588uHPnTtM0AHZyevroydNffPHlu9evTo5Pz1edp+wTIYHH+qsBAbOufd/u+FWvB4DAAOSTkSXnwv3E60T40rRSNXBY+LJxFQg0TO/5TKQvndl6N5YVKhOTM+KeYay6YVtHKxFKpb7oZO5xMLiPdumtG1TczFjWsSAjEgCZRcCAgADkCB21ZAOxR29QRPR0jkA+LUmE5pkv6D82yg8odSyOBoCGYJozmoZAKmJmgRkVTJT9sYOAhdpLM2vmB/OD+QESZzM1EAyvjt9lnnUA8VdPnh8c/PlisWdgVVVVVVVVVb2nagRHVVVVVVXVt6D/+B/+7//V3/rOm4d/+vnzv2ocOIajm0cHN45Aes0p55Rzkiw555QLkF52XUpJRMBYxbJoCGwAktWVUi4MN6GqZhHPrMg5leJYSCIiOcfYEDEapJQkC5i5LZqYxbTPYgpMoWlnyUwAbxJ/ehRJD/qzhWU56aQHyDABCUU7PlkEFVERdMIbIzENZf8YFVUAhvgNmxzB1Ay1EC0z8whmByCo/ppjGdU1ZFTVnDMiqnL50gG0JztnATNiMjUDcyf1wHQQAFRUVR1JIBabH3tQteMShX0SRDSArkdVRYDUN7O2bdu2aRpqW9E5IHMIqevL/cxpvXD+ctlA0GzCZ9DG19+LsSKgDRDbhpX2Qwf7FnsKu32Aj3g83XU2uv7h1gNuks2ygVk3LsSGAfON/BNXYVzbGLgXxV8UQHhJFrSVqYUPaaHicDu/Dea8efBLe2AkxbiGnhMz7rfYiqEDh2GF105WmbYCN27QBNX6ixuO5j27r4c0wlDvb+oBB0OEZsZt28zn83t3737yycPPP//8wYOHR0dHOeXj4+PXb948ff7iy68f/fKrr0AyGBhFiszICGaimkXV/J2KXsFP1Lz+oDnlBgDxcqrDM0GtvLs3S5v61qWrEEve8vrJo7guvmpWjrM72WIA63cT7Ju42u1y0wFACziABhizQHAjSGV9wskTw9DpM1BAZDMGKNHPZaQD+bIeRCTPYsKGKCIyIBNxmbEyU8+gAjNQR+PoT3SFwZAvOZOpAnsvkAETMXIbOAQKgRGMyGLA+bydz+fz+RyJkkFn+Ob4jJo2C2RewYObD56f/PllXVNVVVVVVVV1XVUAXVVVVVVV9e3o/Paj+ere1w/+6Hde/lsnXc/HJw9m84PZQWjzDHS0bpmBiohKFlUTydKvct+nlIRDMICcJOecUur6Pqecc+66PmcRMyIUlb7ryjrmATQgoBqoCCFacDKgqtJ1fRbJaiqKBv3qLGXtRTs0xXiE9OmtFkS1XywMOoA88KcLSZPKYGkGD91o29ZrdIUQCFFVc9acpdQoRPS2ZV8ZjkiETAERU85mxhN/Hk4Y7oi9vLahc4kQgruYvYajR6TGGAfcUmKXmbjES4fgmaqO47OIp24bDj23g+JUVURiCMXyjGhqItZ1vYjMtCUiAzg4mN84PETA88Xi7PT05Phd1rTba3u6cU3McGO7D2LQI7EaPI2wlVkBmwkM1yGP7yUc0NXaVQ2o1ziYmXkFtitwsAoAAIfCy0QKrHqPFhJMTMSXtGf8bHPqZON0m5ERVxLZDwXlomYKhICef7s5qfBNNFLJDdI60ZrZXm9C5YMaAZPeRsJh2MP+Jl15KH+q+mMIhzs4zNFtbz/Fo7bhDjbTYuMtzVBA48B3bt/6+MH9hw8/+cH3f3D//seHhze6Lr17e/zkydOvv/760eMnr9++W6beEJuDG0RBszGTP4XQAFRzSoZIgbNIFsmQ1OsNEnhV0/LwKpH6znnNEAF4PYpw+DgEbqhP3eHggC7PZTEzJAYzUwGi7ffLkP68/oj7umraZ+ADXsHUoz2cbF8+aTBZ4mFYatpCQAzDx+hGZ0RAIKR2Fr3zS43HLMaqiKCoAAkAQNFjjdAQEG20Qw89gObVfUGzx9U7bGeylqkNzdGNg8MbBzcODwJTE7ltA5qCGUfuRRddfvfubCGiHFIWSDEfwR89v/gKq6qqqqqqqt5H38iWl2rUAAAgAElEQVRCUlVVVVVVVTXVH/4h/KD7V77b3n/9jtv5jSa2N24cHd24ETCTdIzGhETIzAiQVYr5LYmbtxRMVUWG0n8ioqKiWQr2FRXJklLvtKHvk8NKURORnMS9aCqSck45pZRUVQFUCtTIor1or5aAe6OzTk9W8m4pz45PX5wuX5+nDKYAAsVkZ1OrouO8MfUVEZA4EIfgxRKZ2T2bow3RSnI0AKIW+2/x/w6OZ/AaisSMhb4YAiB5sgYWz6CVQoJEVE4xlBDEAYO6ow+suOeISMRZjB8Mc87oB8bSvV7aChHVVM3KYnnVYupGssGZTYRu9TYzyTJr27ZpYmxUJOWU+m61XK2Wy8VikVKnXo0SJqDHl5YTrf2aWP5vGzbNQmyu6zXeqjC3CU6nG051HZTpVtBiR3SDsiluNBVg7PmB5A+oVM2HStlTnQJvtXLNrNcJGzrU6RwP44OvQFhQ9R3WF7Z2Xe5xto6ntukgvvSy1wB65LB7Qoen9HbfvbKLdrxaiAha3iuG24eappG875GHlpcxubdlk6vac9EwvKEn58a9n+7Zcf95AEoKPl61hmDvuN66WVgA9JiKDGsOCj6kTMCTK9QQiIAQGModFS+ChwixCYeH83sf3X3w4P5n33l49+7dmzePmjjru/T27btnz1++evX67bvj05PTs7NFSpJUBSzGiEg5CyEiIRODqomqZgNAIkNUNc3iPmXAyWNiuC8Oof3pWlYwmKI/92BoKRgSAZKZAAAQlQFJJVwDkQHcFDyM49GlvKbuE8uy+puspCQNe8CwOsFUs6mAhxp5D2/fkXGqq1zU8EMCAlFAYsCAxEgMxmZswEDkDxh/bhSO7FDb0IwQCICG+TgET6BWL0iIZojETDEwooJpIAzETQgIEhjapomRmhjms1kbYvApAUIgVBVQIVRCRGIMgdr5u8Xy9WJ5mmV53r84lRjwjx8/u3hAVlVVVVVVVb2fqgO6qqqqqqrqW9Mf/iH8iz+8v1hh23JKy0XK71bd0enp0Y0blDvMq0AWIzcxEJGoMBMzgxoThxBFRQEYkTkwMXhgshoiIBIip5QkZ3FbmNpy2TmHzSIp5ZRy4AiAknOfUp9SzslNdSomIur50ApZqRfrst5O1ht1QHdetTdeHTOen3b9IgsMkdCTzAxPzhzRVaHAniISgphGi8ZEyIGIYBJlioQc2IaCV75EnD362cxpb4gR1GxkzUxMjAMp9kwPT2QmCu5TDiEgoooSEdK6YJ1DZ44MGQGAmQFM1dgvBNFTONSM3ZCNmFXBg7aRgApLRUQCMjTRbGoKliWpqINsADTDGMLB/DDeutmturPT0xDDarlIfZdVVAaaPvQeDpx0XGlfiO0W1b1uyMRAfDZB0LdiLsAp3C2k3OnVVTti8aRON9xyYAJ423Gy14C9EHzqwXz2YgB0xQ9KuL0XDih2m4aNRLIg8mv1y+j9hQHB7ieiuN5o763Cnfa8l8aqcWYAOtpUL8qGfh+VGzug2d1vr2MZdu8berTO3mFwuRV22ym78aVd3J7pVvvPWB5IflUT6G8b/8AwxkylEG8zMg/nGa8HQ4hNG+cHsxtHh7fv3Pze9z7//LvfuX//o9g0kvX1q7dPHj/94osvHz999ubN277PXuiVmRlJJUsvACIiAoCEEtgjOMzE3zsUAgB58gahm3RH9+4waP0FYvSCemamhkyAVN4TZgCKxEikogaIxKVDaAriAcDGWaDxDtg4qMf+VgMxnwUkoiGaQ0GHmA6fCjItUyM29vieqQhEt5YD+jodhBYpMrPRkP7sWNnfXcPb1yzl5PNxXl2WEERNDXz9C5Gn/fvwQ0QkAyaMgecxEhqhRqImcBtCDNgEats4m8VZ28zaWWAmhL7rV3236nr/4WiSm7aN88M+dWnZnZutjHLKbxcwj7RM+xOaqqqqqqqqqj5M38ofKVVVVVVVVVUb+u//9r8LKcQlHx+KAphAACPtsTtrIzGaL4xumjbGaKKM1MTYti0xm1oIITADodfrAwSiEGP0HAsA8yqFqp4wYSnlnHNK0razwME8elTFM5RTyqqmg5C4nR2eL7uTk/OTs/NlL51ij/x22X/56u3PH738+uXJ0ooJWgFsbfccmVSxuBmQgTge8KKHHNhN0YWWYfHcUWBRFVME8GpSpUFmiG4uZhXRLGOqg/NlEQGHGoMNVrXEnJY2TVIgpgEUNnBkJlJV70j/FhMBQBahwVedVbKIp48ykpaUAg8s0FzICBGT43IHhKoWY5zPZrfv3GIiyTkESimdn50dn5ycny9yFhUx08F46HQWEQCHXJECn0Zf+XBRV46x0Sv4vromuCzwq+Rke8WzjV133bglwrW4Nm13y/IlwWBhdHflYKCGdWk1M1UpkQTjfuUUI58dzl4SYTdOwSOiLR7tayLhbwKOvyVtZm5YIb6I0++6PswHjR96jXZBaDrAe9Pj99f01Fg6ZBtrD3jdjIYnlz8HSitUTTMxIzEDueNZ1xMOeveju9//wfd+8MMffPzx/diEW7duzmbN63dvXr589fzZi6++evzq5evz04UaiIFmI2IkFlFfjiCSAczTe4iJmP0J7KXwAMAJLw9v/vE5M70yNfDSrOw42CP1y3KPIdVo+EeymD9RBziLhACWsvgKBh6SqL1/iEnNxEpGv3n8hxmoMfqyD1TzAKeski2LmpiW8oNgCjvTSwOGHt+VHriBjByQAmAg9BqLZEZgYEBmkzkWf1LYuEoC0aiMUkMERuJS0wBDoBi4CSEyBaaAFIgbpoY5BmoCB8ZAEJgYwTS1TWDCrluBGSJIliySJSMHioEDH9y8hcwv3p0sxFaGy7w67pbax/MF/PGTJx86Vquqqqqqqqr2qALoqqqqqqqqX4v+yR/89RNenMk7CneSaE4pWooAsDpDS2Tu2/VMDgxEgbiZtUQkWUJgItISXhzUFInYqS4WekHIzAEAHRe4VzqGSBQG75+BgTjm1eJHNlUibmfzLuXFYnW+WHUp9wrK8Szpi9Ozr18eP3p1/OL4/M3p8t2iSwACMLHMjfCKhi+10EQiZi41njiQ29gchwC4h9nAcBSgmToZIURi9pwQcnuy6hD9PJ7aLwq0VMOydRIDFge080pTAwRjcJ4CjnDMENE7yiNQRBVLPgfmUuMRmYiJxjJeLpFMiMw8xncwonN/RowxHB4exBiZ+fDwIAQWyV3X932fU14ul8vFous6KRBqcEAX0jqaoTeqjeEuXJtosH6iXYNT7+qa1JLKJIFPACBxGBH/Rju32oY41gu8eJvJRUD53ONXhrwU96qWtIG1y9j251qs0xs2zoUTz/YwobC16zXB6La9+np7Xf/4W4efAOjJ8B+d4Fv24fc+x4cB6MFnfgHJ/7UD6OkhRgC9aTV3E7EZegRHiXAZfMbF0D4Y7Q1BjRCbtrl9+9bdj+7eunnz3v2PPnn44Nad2zE2y9VitVqdnJ48fvr01avX7968ffPuZLXqUREpGJCqEjEhZ59kQlBTRAgheI4HcVBTGekzkRkQYSAmIiwrQra7Rs1EtCQ1IYKBliQNnMrvvGqZevFJMZ+um3YWjpErw9c63ML19JWaqbKbjBFUxSvNmoipmMowD2S4L7xlmCfB4cZ4gQKMyMEngsDQSye65dzKww4neyMAg7eAoncrIRMF8jmpMjMVA7cxNCE0McTIHu4RkAMho+foi6lK7sGUmTx3I6UOzYgA1GdAkZqWZzOeH2aD09VyKXaec9fJuZ2jYSfykz97+X7Ds6qqqqqqquoqVQBdVVVVVVX169I/+IO/gjTLRr0pZs1dptxT6tgy5J6QUp9FJMbATATEzGqWUxpoQm7btm1nYqoGiMDE5BgUgIhn7RyJYMxHZoaSvlvctcM/VPI8B0NoCMG8NmDWrJrVkuJKYSFy2ufXZ8svnrz8xaNXv3z67kw0FeyIAKDDMvC1321S0goRkZlD4BjY3cJERKSqXdcDOewtpDiGAADZY5oBmMlNqm5YzpJNjQhDjG4DnyQtoKqJiBNqVWUmJHKTa2ElBMAYmH2D8Y6oqqiOYBo97QNRRLOI1zYMDqCH/vLV6MwcQgAAEen7PoaABiklM3VbaAhhNpvdvHl0eHjQztq2aZhZRU6OT969e3dyctKtVpLzxO6LUMqveQduOqDpwt/QcB2jjTbches4pke9lwN6ANDk1Rf37js1oQMAbsHCfW0rSSk+PLmMCs/OHgH04L0GGpytOviYx5FcjjaNWUAADz13VmtlyT58KIDGfZtdx3u+d8fraOvqtizPu2T/fRn0LoB+Dyv9FUnNF+313ntcKgTwt/BAV3HyHQPPuHASvd6nPCdRTcCMEAPzrG1v37r1Wz/8/m//7o8+++w7RzdvENPb45M3b96+ePHy68ePHj1+8uLlq9VypSIYYgxNE2dZTEQdQCOSqKiqh3sQE4eSPk+By/1C9HwLFQUA9icXYCHLOzMKDqD9p4CpTTej4aE+ziuCmpoFZjBLKfsamdiUgn6SM6Ax83Bk8YQLmNx0M7Os6xOKaM7F9ewJMGZbT6jxE9v8hAAIiAEZMDp9JgI1M8WyCsEIjMqPECRf0uA7IgSiyDyLTRNDDDQLITIjOrlWMI1MTQwxcAwco9vJMRiDgYqspE85Sc6LxZmpzucHIVBgZ9nAZGTWhjCftRBbmM/PunzSpw4xiy2W/f/wJ7/4V79376Nb4Z/+Sa08WFVVVVVV9e2rAuiqqqqqqqpfr/7eH/xVysIqnQCB3jA7OGgDoObUrbrU90weSkHJozREnN1CwXAKSKKWVQIzESOhigJYCEHVRHQ0IJuIZzyMNrkhOnZNNIkoNI07pgGQOHBokkEGFMTeYGW4Evzq2fHPvnrx+NW7t2eLRZ8SgAAKlhXYOECeCYBWcIMz+8JoZo+4LtC5uGJlQBaB2cxSTqbmxkAaCLU3POcEAIGDm7gBzJM6sJivYXBPD4W3Bl5sZoiAjM5MJeeRg0uWLNkXwiMAIzvQ8WqPG9R+vLTiqS6/M6mZiBCWoofuwkwphRDatg3ByzDafD6bz9rZbEaIpiYiq9XqfHF+fn7edaucsg5VyEZz60QISHCBRlO4FW5TXrz+gLwurzRzZ3vZx2xfU8HMfAIAvFyk+GL/yZam6yqC+1oyXpCplfkS/0LVEdYYjTulz2tNazYO/6oaAhCjB7ZcAvSv0Q+Au8j7Gvtd85SX3w5npmWSQod4meHjxQz6Ep8yXuKAnu42NeGvCfWvG0BfOThxYp+F8tgpn27dHC9n6nM8ZqbiD6gmxIP5/NatW9/57NOHnzy4e/fOR/c/un33dsry9vjd02dPnz599vLl6+Pjk8Vy1fVJzA3BGkIkYgQUMVEf+YGZxMTGN4gVXkyERGy2xsc03EgryRv788MHZA3+XFIRFSX2AJ+yAQ5FXAHAVEGEQgAk3ZycsDKNs14pUWYScfP9YsW2jB7XIWJZfEeAPfR5425MPicAAmwgMBACEBjiEEc95smUtR4GAAGRiUMIgYkJGSkwReI2hMgcmCJBQCBE9hUjaF5B0MshesVeE/UoFTNTUCSkQLNZG2MAQAQlhBj9FIAA89ns9q1bHdC7xfI45WS0spxzennaPTte/MXzt1cMv6qqqqqqqqoPVQXQVVVVVVVVv3b91//hv5YzmFBoJRLems3uHh01bdsvztNq5UCTQ+j73mv6FSsnUd/3fd8jclltPZA4ydlDKrJoToJUlmRjySHYttQNKAbd0BqadgNAc8xgCqAAGVCIKc7fnvbPXp09fXPy8vjs1dnipM+LrBlRoWQZT0rrjVjKT0+ARMWsTQVDDwEONqwk96gNEVH1anPIgZnZoGySJZv5unUd17AzFRYBCCJiBiEwFOuzDYzSrARU+EJ8c6AvIl6JkZidcjIQIwGgp3qM1IZgnblq7g8cUjmGTi1d7FXxcs5+B0XEo6ZjDG3bzGaztmmaGIko57zquq7rUkqqmlPKOUmWlFPKaZO7FRw0dOx4Qhz/K5vhNoC+Fly+Jn/2GzFOhAw5ADtHMhoKhJkMmbprbFzA3HakSCHU63vmh9vsdiUcg2FLlPPey1ybhceGFduph664o3zLmT2MFNjadfOFEthwgfV796WNnvkWVKZE/JhmNpLHARWPLu+Ncxpc3IS9UwG7n+3er6ERu0fGC7/YOf5FWlPjCzYYmSlP7o2BiX+FhcmPfNymUxMIGBgPDuY3b968d+fuvbt37927+/HHH9++dRMADSyl/OLV66fPnz1++vT1q9enp2ddn6xkzwQojxFGRPPifApmwMzkABrWI1NEEMEDiMDMV2D4fSRkQCjp9zA+C9cXPR4HAb14rKmoKDKNT6dxqq3sZgpqGAIyFdRu09upiF7wsLwtfaHIOMHmBy0+cjP1zA1PfIZ1aMmu5Xl80blzACzGZ2ACWv84ACMfwkN0tWN4BCghGyEWkzI6hsaAJXkDVQmM3WdOQOahTZlQvSKih4SQlkwWDhQjxyYeHs5jE8x97oHaWevrhqhpQ9MGplfHpyeqS7OcoacTlGiCP/7jX145TKuqqqqqqqo+WBVAV1VVVVVV/b+hv/fv/+sUlBAx4J3D+af3bj+4dycQpeVicb5ExNg0qpazSJaUs9eJ6rqu6zoAT3zmru9yzmbmnBqZcv5/2HuXVlu2LL9vvGbEWms/zuvmrXxVIcqyGgbbmAIZIzWq4a+QbrghhDEFsv0h6kMYgRpCWCDJVDYMdqOaFgZbWJAI2aaQTKmUVXXzPs/Zz/WIiDnHGG6MGbFi7b3POTszy5m3UPzz3p1rrxUrYs6YEZE7f/M//0OHoaSUVLXvunB6QZjs3CFCJ9RMK8Ht+05VObXgaOalmLmrgYEV01xKMTMHIEFuidedyttt96fvrn52vbvaDz2AIfo81wIr9XjU46ArxCycJDUp1p1HZS1EROQZAUQiJGZimgoMzqMGThIekONXVUWoSakPmLu5FiswFjzEiWlOGdCI5g4WmBqnYAszm3JUQx5QpgZoGwBMXagu5jiimZkNORNi0yRVNVNETCJNSogoIimltm2bJomkvu8Ph8N+v7+7u72/vwXzI1GKPjMDoqtWaycK0MNuznA4Bm33ctL4p/VUjPJTmz1yYT/T/YoED5j4z/PF+XePn5zU5XsCByMAONBTcBUAnPDxbqcB/QWP+MEOPT/U4nGr5u88gd19fuvVD549qxBbPj2yOBbI/NAOwOc3u498d96hJxD3R1v3gfKGdYMp82eak6gBEUE0ySEssVFWL3z3gADjPXtxcf5bv/WDv/bX/v2/+lf/vR98//svX7zo+3xzc/vTn/7pn//55z/77IvPv/zy9vb+0PfujkScUj3yCXKvM3ngYAZEBAThgIbTa+Y4KeDjrGB9Do21N93BPaboRqQ8zi0ce+11DyO7nR5TEb4BHvCVSRgJEcmKmhnVeB9wN2JMKdl4uKn0K1QgDWCqOXuspnGvxQYBEBwfR1Sf/ooACbABbIETkECthzhetO5gwomZiYCZKNKmEBkpQuyJCMEJgYAQHMHQParfliG7WRJhRARzLSXn3OfNJrVNakQInQlXQo1QYm6b1CZpUkJwZBCm1bpdbVar1cYB1Zyb1c399u1ut3frSlEfuh/8G3r7G9alH/+zzz52jS5atGjRokWLfiktAHrRokWLFi36Fem//1t/XYhbaOnMz9fNy/Pz737nzUoSlMyIEiHI5gCg5gaOALnkPJRp1XQJbxri0Pe5lADQfZ+thpB6SokQi2rOOeehFK2QtOY249Dnoook4BB5CWauDjlnNYUx8tMAS7ZcIJtsC1z35Zv7/qvb3ZfXt/tsg4OCq0NY+wCe5G3hSwyzMxOTSJKURARrBgBW2ovERCJSS/zBMeh2zmumXwEiV8Eq4SZ6CMUAzM1cK04jmn0XIJIiAsgD4WSdjO+e+gfjraIZaqVEAkCL+GkicA8YPdUZC7cvYRTrciIcLauV8V1eXm7WaxGJN5k559x1+7vb+8NhP/SDavagolhjVQADB5GPluL4cGpwPd3vHYjH+lCFw4cj+FD+4PuP/LBHw/K8ec9gkLN9PsmX4ehwf6pRx4O+Z99TvcfZpfKE3/fJ9r8n0eIDfXrmn9ijCfXpDx+fwyPNxxmK/ah9GGYbhP/VT1s5XzzxQQB9Crv/wgB0PcPv3+4EQMNofzZwo+qwjfSIEjNi6NCs2ouLy+9+99NXr16/fPHi4vzszSdvPv30O+Ceh2G33799++7rr775/Iuvbq5v7u93h64UdXBUUwMnJjcFMBJxd1cFiKUdMk5IORIh0fQ8QbdKi6kW0zx5dhG5WQ3BmJ+sMR+mPqzoZJnDZHpGQBaeLgl3x0jCJgRAxyglWJ+KNgJ9d0WiJBKeax4nLdyqD7sGWZQcrmcPa3e9zWfJK6cv4mEaxufk2AA1SALEdQ4IAeoqDgSolV7rQxgQfdyz1ysockIcEZzQCZD8OKXUpEaYGAHcEJwRm4YbSU0SRhCGtXCTpE28WbWrplk1ycGYqVm1DqZu2UCRhwL7YbjLQ1/KLpdshOs7b+/L5fWPf/zR63PRokWLFi1a9MtKft0NWLRo0aJFi/5d0X/3D//5P/jbv2sJhyxNk2+7jr65evPmzdl64/1BhyFSkCGQBCIiJiZvWhijgrWmi9a0aGJS9VxKKcXMEVGSIGIpJdI8qqE5/G6IAJDrtrFu21Urhh6GwcyICcDNVc26rj8chuJyBvIK05vL8vp8vWZ/tz3cdmWXtR9de0/1dSRc7u6gZqpUNzRHJkB0B4vSf4DGVNNJJzLxfgDtjmpWSmGKfGkcPbZVVkGdnaAeRMJaZisqHxIGCYGJz8N7umOmCI6E7AIOarX+4bhjdA+uVAMrbAwaAUBVLVoQ0VTVCrOYGgsTUZKUUnN21m42ZyLNfr8Zhpz7Q859KUVNzR25Zkd4JAVMC9vdcebBHTMiEN8fHj07E8+Cow/R9vFQx2wDB8APQs/Zd59renCYWYCP3GvMAUB4glI+C3geB3luHX9vMx6g8/mGT2Dr9+iXc3q8N1AlWO0jaP7Mw9Uh9Bn+PuYRP4WPT7/75OTAL+1picv5PXuZN7Ved+NMWUzVWeRYGCKs2rTerDabzYsXL7/z6ae/9Vu/9fr164vzi6aJ2S/68osvv/zyy6+++uqbb96+e3d9e3s/DNnMABNREhEDjJnA+tQhGotxAiEg4xg0Y4AIGGk/x4dXTLohESHa6LKPh08xB7CR38Y00vHhVh9wiFNi/4Sb4/E+PXYqgEZkrqZoNTdXd49nCyiMedBxZryu4UCP+ofuVlfHqLmpm9a5jZMMk4fceWoVATKiACYgAUyAjMRAY/jG8apARACPTPY6bQCGADQOIjq4G4IjIGMNy45VLUIkIk0jSVgIASwxt400KTUptSKILugr4SZJI9wmEWEmdEdkQqJhyIc8FJCCeL/f71TVfTC4HtZrHvhw+U/+6Z/9khfuokWLFi1atOiZWhzQixYtWrRo0a9Uf+/3/nPhvuj+1dknyIhAZyKNF99erddrYpmKChJhahpJiYmZJdyyDiAp5o/DEEcIiMLuXkpBOvrpghGGz41ZAMDMzV3VhlxKCd+bFbViYyA0gFlRzUPO/ZD7vhiQOTtyp3B7yF9e3X329vrP3938+bv93aDDVALs8R8Uk2Ox0iOqZmiSlJI0CUaw4jUjlcIXh9U1d+QsUTAQACKcAxFNvZQS7mMAwCeyKdymxeIzjBcYyNwRgJnLoFoUEYniX3Q7xjLUs0iYpOYg55wBUJIwEQCoGUfINREgmMdyfyCCamY3Uzd3EBEEN4/fPJJDRKRp0tnm7HyzYRERSZJ2++1ud3+3vd8fdofDQUt290hHGHs2Zb8iTKv6I1EEEJA/egX+cgA63jqi2583m+I57YkMD3iYfuDTj4/KpkkLgLDVn9pO53s81VPM95mO8f+/NSY0zFp4alhG+BBSn0TTGE2c/wgbP/L1BwsEnrj3n8wDedaoPbyL39eA0fus02TTOEvjxPS9733yW7/5g9/+7d/+/g9/8zvf+fRsc7Y/dPf3293+8Pbt1RdffPn551+8/ebt3e3tuD6kxlsUc0BklvAzi3BUtpOGzbTkDADELEm0FC3m4JEa5GaIyBz4FGPKzc2FeXqeRE56VB+l+sRBQDC1Usp0F8dpgDHWe3qyBW6OUGmH0X+NyEQI6O5qZmDgwCLEZKWuyTAriECCprVAKE6zCFOu/dH17McX7xk4RGCkBCwVQCM7UricHRHAI1G/zgqOHuejV94RPNKfKQoSIhA4IybmRJyYG5bI7BACER4BNIFbEm6bdLberFZtm8Q0o2nDLESEkEvuhm7fHcxczYtbl3tDSetNxlSIlCGX7vDD/xff/pXD3Zv/5Sc/ec51uWjRokWLFi36C9G34u/pRYsWLVq06N8p/b3f+x09/ytfX/6Hv/32/xAYtHjruhZmV9TsrhNGkpRS24BXOhGLvlPTBARiZiRGJDWryQh1UX64b48MN6WEUJeKu0NRs1j0DOgVbsZKaHMr5mruueiQFYnB0Qz64odBb7v8bnv4+m7/Z+/uPnt388W7m32BwUYMPecVJyZWHN8iRGZmFgIAYk6pCVufO8TybwBAQqDwFoLXteRT1AAiYLj3YOL0kztylGN1QMMUtxr+wYAv9fSgF3cLe/hoNjS3J+JoHdARQLWypHpoxFjFzkSAkaBLAK5mUUNrdAdjkJ3wIUbH3Q0BRNKqbVftiqNOIhIROpqaqqlqycMwDEM/5K7raoFK1cq5IRbBh+0ax5M/najjSDzozEdjFmbdfkSHfTzICbt8cLCndv4+M+9TcHtOUacE3ec0+PitORh/z1fruI8fH33w0zdxdAdPX6GfrxnPaOh7Xc5Pb/sE3p1u+JM5g/eeMQd8lCjyeGN/z4A98e7xSvDZRu9P5EwAACAASURBVKfbPcslj4/eOskgHldchGnYACxK5F1enL+4vLw4O7u4OL98cfHJm1evXr28fPmyadcOuNvv3769evv23XZ7uL29v76+PXSHvh+0aI2br1XxQOORQmxBokXMzd2JMeKlo2HEZFqrCDJzJDjP2owIaO7gQHXO7+iAjiNOfau9Mh9t6PUc2niiI7pi7oOOpxfFQgcfq68en/80fwA4uFsBBCbUohYpIuMMlvt8pE5fHIfyOMjjRCIkpIScouqgY8xnTOVoI516luNRneGI9bmOGOUHkQmFaPoniTQsrcgqpUYkCbspIqTEQsiIboroTJSEExEjmBbXgmYRfqJg6q7u6rFiRWSzMaDtodNGFLjrM18ebLUrl++W2I1FixYtWrToV6wFQC9atGjRokW/Bv3+7//+q/2fb/qrs8N1r8VNG7d1SqADlA7B3U3VWERSMnVzc1AEZJGmbVXNzANAG0AeMiBKShgkAABmaAsRkzSIGJgCAMakYiZmIkZiQnYA01JXQxOpeVETEQCwYv2gg9rg1DttB/3q7u6PP/vyX/30Z1d7v+u1U1WPNdUAD3yRPtFKRKiAJNBsapr1epOaRCwRrBGwBgmRw0CNALF0vIJpwrrO3R3MDQCFZcyArjQx2Isfa31VAM0cOaKOhA7gZoQcKOd0U5/vyNxKyQgQeBjCVO6OSE1KOech57HUIYmIuQ85CzEzM1VUVHIO2zUgEGFKKWgyMzMxj0v1zez8/Gxztkpt07YNs6iWrusPh/12u+u6Q8lFh8FKNjXzkTgjAo4r3wEf1XN7HKrw4ZiFiSGf5ABATAZMAPpDelRLcPQjf+iL/sSrucP3CaP0BwI0Ph6HHLG8x12MPG4esDG5zo/bP6cDP5dcn4WgcTyLj+OoJ2Q/A9AfdG37U589mGj4BfozQ/gnDPrpHcWsDGBkOp+O+SmAnp5adZ6LCJmYGYU5Jfned3/j+9/7jU9ev/7kkzdvPnndpEbN9113fXP37ur6y6++/vrrb66urg+HYRi0qDVtE4RTVVUVZ+VJw68bjmoSHpMufCxseDxR8ZGMALpS8UqiGcfgiXhWAAAiMk6QdrqRAMdJjZiBC0038Fg/tc6NlVIAIdJ7AMDNVM3NzJ3isSlsGkUIuZJmL+hASKUUKwrgYAZjodd6YJws8fNROy44mD/BBSqAFkB2IIjpuXGMgqLHMI3AOrgzETOhEDJzLNQR4SScRBJRpJ8kloalTakRTsI5D26FiRgBweN/ntzcrYApuYEpWAFVMHUwSkIpcWqBmJuWm40R7XPuwHPR2xWuM2L2//Ff/OtnXtGLFi1atGjRor9ALQB60aJFixYt+rXpH//e73agHXvKxTKswFshygNQASil5PCKmToAIGPOAyCkZlVyKaosyQHNDIiJiIkChMyZGhGJiBZzAK4WPIsgCwRUc4CIFmVwUNOoB0VEBqAOwoIIbp6LFnUFBBZD3ud8teu+vj189m7/+dX2y+vbvfpg7ohRn3BGLcK2LFihpkH9B4mIhFmEpUmpdaSJmAOhu4UPcSI7UI2+CD6msCLQWASsBoeOFr4JCBGi1zXhXpFjxGGYiQgROYCZqpq5ISAxCUusjgcAdyu5EKGMiR8Tx0fEKWKbmFmk7lmLAxBSincc1NStNgkBmFkrJ6LgVDGjAOAiQkyIsFq1q9VKhJOISOIxIWS3227vt9vttuu7YeiDvEd9M3CP0oiTJROR3MyRgLgiP9U6ERCn85hkfTzBODNjju/BOJSP3zyVw5S+MgfEDw7zxNeOvGtuen3P5h/TRx3TcaBxnmH0i8KEvP3Y5Of5r58iw89rKnw8tGRMCp6btR9g+tjVlNTygTOH9SZ60IjHB31M/OExTZ7f5j42zAHsw2ejLuioqBS91vHzcVoAa3dg3FuEOSAk5ovzi0++88mLF5dvXr/6jU8/ffny5fn5WSJxt2EY3l1ff/XNuy++/ubq5vbu7v6w2/VZa/C9g9c0DMIxXH5MM/fTK/64XsJdI9JZiwI4MQEiOMQEEhGZ1gh4cI+Sq8eAmgk0H//LJ/8xhDN6ym2fQPz4Do2nYho5NQMHZgYAcC+qDk7jxEg85wCciKPKLFTLM1hRVR1zn/XhUI+FKY8p86djTAAJURARgB0YsPJlr2ZsHGca6xMWgMCjnmKTuEkiLMKcmOIRRwQpJWGRMYuDEGMhiUeAkelQBi0ZrcQ6HTcjJCLRMhDaKnEjuEp8tmoTMws265Uh9kXb1Vlan+264fpwOJh3pRyIGHxI8D//7wt9XrRo0aJFi349WgD0okWLFi1a9OvU3/07fxN7846aVBB9w3K5ltVmA5i1DGiATtPi5yH37p6aJmctqkiiRYsWlgaJwEFLMbUZgHYmJua+G8LrV9exB4c2rw49dyIBQHcz01h4jsjIXBd3u4dBr6gRCwmrw6HYfW9f3g5f3h6+vN19c7e7PfTFcQDPowXaI/ECiEAAAsZOAHqKe2ZikdRIalgSTPUSwzXMDDgjgMGSK67CcCXX5fDEsZmqAVQUO51nr7UEkZghzINWiwGO/Nei/B0RMTEAqGns0IrieKzqRqwmb4R6Sj3Kjh3BtzsShX98Zq32OCMYyQIeVnCrJQzh6GM106ZJbdMwc9M0bdM0TRPB0+5eig5DX0ouJfdd1w9DznkYBisFptGq6/cpzhOS1GpktRxY2JynK+UhK55qo83ei/H8OCutBcZmOz2FaE/88fk+XvohjvpLa9z5KTh+gpk/avBTrZpXNvy5mkHP+Mroi8XRQQtP+4pxzHX4CA3/eKVKwEcW6id909XnCpEofKwAGj8fnczpF0QGMNNCQR2nG2RMQ3Z3RCCAlDg13LbN2dnm4uLi8vz85YuXr16/Xm/Wm/V6s16rWs556Pv7u/vrm+t3V9fvru+u7u53+0Pf96Y2RgxNwUTTvIOf9LSuosDJ9hs/zS0KmAa3JSZEAsB4ohKhFXVAJD7urB7l1NVfT4g/uNyOg3GcSIiLYrLc1+cDIpqDg1Nd94CmBRyQeETluX4fycHMDaM74ZOe/XM6HMeoE4cHH9UxJoCWqCFCB/LI3KjW5npywXGsixjwnhEJkRHD5syIQsSxjoTAEYSZEdEBTN2MEd1isUtMRbhZBjdBJAByBAQmYUkEIAyrhtYNrxvZtE2bEiceTI0IOEm72e276323d+jLMFgB5EL8P/3zf/XEJbxo0aJFixYt+pVoAdCLFi1atGjRr1l/97/8m4lBWIj79ap5c352ebHZnJ8xEaiiuTADgoFlLQAgIkWtqIFBPwxDHji1iKhquR9K1ol7hDkXALtDN+RsOhJVs1JKKQUAVLWUTCSIDACqJZeSh8ySpGn6riuq7p5EAKDveyIK/102OKjfZbod8Hbwn37+9efvbg/F9waHaUV2RT5EHnXlojagHfEZBtRERGpX69V6Qxwo3Pddl0sxMxIm4cmx6EWnGlxExMIB3IgpvlhynCUOBq2m4ak001rIayR6SASIeixGFp9j9UubETMyQWXyDgDENKW+xnkIXjxf1I6IwbIDQMNkKHaPomFmFpRGrVqVRSTeMXNVzaVEecNwSYtwYg7W/fLly/Pz86ZpUhIivLm5ub27vb+73+52fddByUfDOCIgOTIiM3HwN/ePU90xiOB0M4STgXuvAhueAsfnJTg/kUT8iwLoZ37xic2m7IgPJWV/MOHj2RHbdfPntvQ52z1hX31KzwDQ8FQnntj3EUADONSUjAhgn6YrEB8dkVkAXMswC3jx8R6MqR1gwiR8fr65uDh78fLF97733R/+8Ieffvrp+fllSs3QD7v97ub6+osvv/76q6/v7++vrt69e3d16IdiACR1gosYwN1srBA6jo5H8T0A5tF6HIsJOFJ/wGaBMxGubxYebeKEdeFFJB4bICEnRAQzL9mJAAngQRjOzC8+aWoYnEwIjVNEPHPoO7gDMSCCKRIDs5c8dgHBDMpwcrJ9vOkdaneeuopw9C/DDEBPLSUEAiCHFXNLTDZ+6kCEzDTRZwBARBZmIiZkYiFiAgYKwzZ6bObmlk1rnL+q5uKqjOEPByZKiVIjTJ6EV+1akBhRRIiFRdar1Spx4jBBMyM0SZDw69sbatrUru4O/V2fe4Vc/O1N3myAkv34J3/yuO+LFi1atGjRol+ZFgC9aNGiRYsW/fr1D/727xr3hYcXciZts26aTy4vzi/OKWfMw6ptOLEzmRsQEkfUBiRiU1NTblrksLgiOuK0vt69FM25hD86nL6qmiPCw5SJg5+WEhEQaFqyah5yMS/mJeeiqqWYm6nlkqfgXHUYHHaD3fd63+n1Nr/b9l/f7j+/3X51fygAUXYqzMp0/JPD5+bM+goRgIiFWUiEiGONPBIi4VTTKrgUI8NYjwtmVQjHEosBXcKRTOCuqlERUIvC2Hh3txFAT1g2DIPj3lxVWZiJazGxqNuISERxIBtpDiESExJ7BLKCj6kgJyvooa5hR50AtFYneF1TD66qaqZmREyEZkZIwkwU9buQmCO2ZLPZbNabCCohxO1uN/Q9mHaHw/6wPxwOw5C1rrVHjHKFz6CdYVk/2Sy6gKcbvX8HjwH08/VMVP1R/bzk+vS4FaXBmL37sb09yA/5+brw7QXQz9gDwsw7WwH0aIL2Y/DEE8OKlXtaTY04Bnms2vby4uz1mzefvHn95pPXL1++OD8/T0mapuGUcrFDN+x3h5ubm5ub25ub25vrm/v7+2JacsmlOKABWuRXUC3WN1rCj0Hf1XANOEVqAHhE6VS/uR0na8a4DAAAmyVj1MgLjzghjpgPRND6HHrU6ccA2mcjW++zujBkfMvHzcDdImjIzADREawUACChWEwBZrUnbsHcp9ML9t5ZE6yhOcHg61iENZsQBUAAGbAhbpDQZxkudbbgOHxxmuLkECAjEHicFgJgAEZgrItpkpAQMjiYEUKbUhJJEnkdzARtw4nQ1FKSpmmbtkFmB9is2oaJXIUwCa/a1f1uf7vfUbsqAPdD3yn2Rbveb7elSThk/8M//uMn+75o0aJFixYt+pVpAdCLFi1atGjRt0J/7/d+59Vm9Z2X6atvyrpdNyldnp2frdZcegEjIRSCKSkTgJFaTpF5bEzAwpKEEiEfF887lKKlaEoJEaPoVtGSi4Zpt+afBiIwgJpHrMU8F1Mzd1e1+sVSVDUyPNzdHBS8y9pl3Q+2z3R30K9udv/265uffnN9vdsfclGH8AbjjI3NKcjMNIwePJkFmSK/IqWUmqbGhECwGRISGHFzkGYidIdoWwDicQl/BdNhqzSrwdNQbcsGiAGTYMz2gMpP0N1VNeI4IrrkCLij5fEOjHmxTEjk42ZRfmyikWOuQLivoS71H13GNXOgZp9WX2X0QlURkIkADBGYuHaT8GyzOd+ciUjbtuv1ehgGUxWmYRi67tBFNMcwlJxLzsOQde7Snkc+z/+7gtfTkZpA2glMf9+F/ASAPoZdfFBTzsfx2yOxG2MNHuwQRg74CxqlnwwJOT0yuPmU+v1h/WLNeA6A9smX/bEN52sL3nfAWV3QX/C8TcZnrDEbPjZzDqDnN/fjlhoARGI5EjRNs16tNut1s1q9uLx48/rV69evX7169eLl5apdsbCWvO+67e5wfXd/fXN/fX13e3u73e4Oh0PXdXnINSKHCIkB0dwj4MFMp7vMTwXxOCAaDdD16QHjUPr4Km5qJoKAv+NdH/shqqEccZ0Q4ZQ4f7xoq5n6wQkfofhpCsx0B87s4bUp8ShzdwB0BC0FAFjGsYjnuJuqmhZXPQLoB0eZvcQpNGfK+gAgAAZkxASQkBgwfqIDHnsx7hp9+h+d0UrtVKMzIKoqMoIgCSJzJexN4lZYCAmdEddN0yRpkrRNSkxMuG6YEYa+J2ZpUrNqgdDMEhOBoxZTA0BpV4es2yED4y6XnqArYNBpL8OA/WALfV60aNGiRYu+DVoA9KJFixYtWvRt0f/6+7+73ZkWGnrgVctAa4YXq3UeeisdCSIhMAA5IwpyQ8LESLjveyBs2hVzQyhHlOdO1TLLZt73/RgkUbHdMAwBSlarlYioWrXAUfUjI/IUyWpmOWerODqwsKm7OirgfoBt53dd+bO3t//mZ1/9qz/56edXd7edAhxTn/2JRemnQiRKDuBmSJSaZr05CyATiBYcEHm2Wh9FeCTD9Z3wME7UOjjRZF4mitwMMzM/xZfVLwkgHBnQBhB0JQBW+KC1lJpkgoGuRje0jTbV+GlmEQYSAbIVlRaNtJAI7SCmGUL10c+NjhAgbBogU0WIooWVqjcptSm5e9O0m82GCJumOd+ctW3TNIJIqjoMw267vbu9vbq66vshhg9p4mITGqxsHCak+yhm4tmoMnb1FID2Dwy+TywL3KvXFGYAGunnAtAfdlI/hZuPt8wTjXv05i+MvJ9ozMf29Gz6DEcAjR84A0cA7R8akQ9rDqCPt7W7QY1vOUlreWQwP9YIFcbVqnn9+uV3v/u973//B9/73vc+efPm5cuXDpBzPhz22/vt/f39drt9d3X97up6e+jv94e77c7UAZCEKRZKjFfChJuZBRBy7mMdwCwwx6Zt4nZ7wKbrXBHVqzBWJKhqxBBFfhEANE0T+0kpRZnW4N9Qp5ROJ2xqu2xa/zFnzw9CmQFoauE4ZnUGKwLj6/IOgKwFwCVyMBxA1WOuMA+lFCvleCs90PGIOI/ggBFACwADJqBEKEgMRO7oTmOTAcDB9VEsD45zUEzMSIzIiMIojIwsxMyYRFLTtEnaJEmYwRmgERFGJmiSNCJtSg0hgpUyZC0KLk0DCO6a+77kwUvuur7rc+eyOr+QVXNQKIIDouKWrUHwf/J//tunu79o0aJFixYt+pVrAdCLFi1atGjRt0t/8N/8rhMWzS2LORIQmhJ66bfoGdGRmYkYmbHWdFJ3IkpN40buCBCZwgwALJKaBgBNLefs7oAQXl03L1rCFL3arFNKCJRLUVViYkksMnr6iJDcPZesqh4LwB0AoKi5AxDnAn3xQ/bb/fDu/vDZN+8+f3vz+fX925vtbTf0DoqoUaqsWlpHhliJWa08hcgOAJEswSzShCeZiOsL5skpDABEWDFa5G6MFkFzC0/36K0G4sghmdgT6oii3EfP5uiphqBCtYSXjh/FQvZqlGaRAFhmVkxVLY5fgz4cVLWiI6rr0rEWIcQRdVUCVksgArJIYKY4ORrJrRNgC42+yyhLyMwppfhVSFLilDilRkSmjoSxPeeh67rD4dB33ZBz33Vd34/nbg6gHXxKyw3S9Kgk3eTpPLLiCaW+L4LjfQkAePLR3AE9c0WfHtqOFtFT0uofwOZT1MPPFfTxFwibnxZ+DC9/9PhHfj4B6A8ebgrQmOU7POMYTGRqZgoQGTccdw2ij+U3bYyBhpMmHQtfAgs2jVxeXlxevnjx4sXFxfmLFxevX79arTepaQlJi/XD0Hf9dru7vr7Zbnf7/b7vhkPf90N2hKHkfdeDOyJLivkqj7AaZh5y9ihgSOTuqhqcHXGcLQKc5lamvOkpRmWMzZ9+VEBs7uGUrisl4ok0ztYBoNrRBTzC59lalJo85PVsn17XU3OOO5gGpDZxakxF5LHqQs0wFm2Ag5nl4qamxVQ9llK871I/LkqIhjpGaEYtOYgy1h4krG8yEsWpqzMiMVkUXwRCipqEwtMLFmIhEiJmSkzCLEQslESSJBESJgZ0UzBFACYUZhGJ0Hpw83huac6m5jGUaqUw4qptzZ2aVYa0LyUzO8mg+ope7Hg78O7H/+yzj17VixYtWrRo0aJfmeTX3YBFixYtWrRo0Yn+i7/7T//R3/mbMmS7uxpev1GFUgprITAwBe0lNQEqKKxwI+IkJHByR3NIksIaLElS27pBmPiO9K0uLddSSs7l0HXMAojhbSYiYkaiUkrwDolPS1ZVcxcWQHKHkhUAmcXMi1opunL+tKH2zeU544ahMSPw20F7qMgiVrDPkdcsEcDddcw+cCtlUKtORWYkQiYBDxJiqu5uhpWfYHVi0kRq7AjWEJEB3CzskEgkLGoa3sPIV0UzAAQmC6JmWj3RRSueCiNz0B4C9OocnK1un6yKAegq6SOsllTCh45EIiKiMdsEIjdAHSf7djReWGjm0xwHME4a5qKMVhwO5UCEItw0TWpS0zTr9Xq93qzXawBXLX3f73a7w26Xc97tdvf396OdHcw9LO1gBg7h5ZxFB+ARkFX74zR+R+72PpCJ048nPsCTj063wulyfQhJ/Ymt3++JHqnZ0Xn6bdETbXlADdHfs13d+Li5P3mOTw/nc8aP9TvPANBQk9wt3PoA6ARgdVLFzcF8zN8I/FrDggkTy6pt27YVkdWqOTtfv3nz5vXrN69fvz4735yfnZ2dn/fDcH+/e3d1ffXu+urq+rDv7u93N9e3XT/kXGqeDYK04u6WC4AjuRGZWSmqasyUWMqQ1azOp8wum2okd4fJTf+EtTzu7tlTA44PTI2Sg+CxqMFAT0/PzMvus7en0378OAr5PXXoKpreq//WnOrpP47MZBQo2wDQo3ppdjNwPXZtnHN5v45PLoqMZkceSTTGczRAMwISg03bAyIGlWZEIWQiIRSmMKUn5sSSpE6UMpEwCSEJMcV6HkdXcPdSVLMVJSIRYeao1OpmZuquCmZuRTOiCUd1ykbWa2lWvVru+p54UDcf/pRe/9Dzb+j5P/rn//qDvV60aNGiRYsW/aq1OKAXLVq0aNGib6P+4Ef/wfe/6v7G//Yn//Bv/WfK5g6b5IIoTKumKXkoORM6goNbznnoh6HPZ+eXKTU5q7m7+ZAHRGROPkK8MJblnJmZWUopUVvPHYtq1/dN07ZtE0g0ZwUANS2lJEmxhr2UrGpN04BDUVN1BBJOqjkPed93iILU9urbrDddvu3s623351c3113ZZTMAQ1A81sSa7LKTrW4kkhP0RCCqVQWZpG2alFJqSs7mRsSE5A5DzmYG7pLSyGrhiFeO2dDxe01xRcQJVOMY+EBE4FC01A3MxvQPHFfXT6o808FtLDs2ugpnebJTMsDcFTlrWEBgn0zFD/5AQ2xECGkcLAcAM1M1HNsTvm8tRYiZw7FuAN607Xq93mw2pkpMm80q2PiqbbXo4XC43d7v9vtD1+ec+37ous5KATdEmo6FdRTGyN/TfI6o5Tj9Nhls6291+/dc6PjeX8YRefQNRJ+CfYkeuMNDI3acIUGHR7TxW6DHCHREeydbPc+F7WAfzDk57v6Jrz44wqN6eQjh6/eT4I64LtzU1FxPpmIQAIEI16v21euXv/mDH/7g+99/+fLFi5cvL15cioiZ9X1/e3u72277Id/c3r59d/XlF1/db7dlKJFgXIoDMZIQiWnWPGBCcIvie4CI0tT4dmJ0wFoy0oHGcxvrGOZdeVwKEBEBZ/0aL9cjpR9P0dz2fzJGON7cxzkmf1z3r7ZkNupPQnAgiNyeGHozSoyEx7ifMRQonpPo5qWAmYNVXzJOh8Z5T44drIfymH9AwMjcEHCCANA+PplrC5lqRVYCIAQCZCJJHMOTmIQprhACJ8KGJYk0SdCrSxpAwQ0RwUxVGQHBw7KtWlwtVrogIwCCOcWjCrFZNc2qTa2s12mzbs7OziQ1QylXd9ub+/1WMTvegzvQgHKL65/85CewaNGiRYsWLfqWaQHQixYtWrRo0bdUDvAv/+Mffv698y++v0aXsI9drlcvLl8yKFpOCQkd3E3dzM2gaVZEnIsG88x5MANEqqum3WNZet/3ENzQPRKdATAXPXQdEjExCQ9D7vohbLDmpkXdjYjMIi4idoiuYRaGUoZScikFSQDl0OfBQSn1RveDvd3u3+76q113u+/3xXqH4qBHxhz9rWxmeg0AozEQa3FAImJOTUqpAahZqIgMDiVWnYOPZQWf+COHpizmmTUyqG5kCsRHYXw21TjilGF8GhRx3EOkT0wfThwZcWJGNi7+f4ibcJ5AMSIte0QlGSuNgsnXjTS6vWcBAmbCzMTgXsqgpazWq9Q0zOLuKcnFxRkRM9O6XQkzAHa5z7kUVUQys77vtBRTzbn0Xdd1h6EfiiqG6zVGDI+O5sDAOGd8TlNP/Ni65xDUR0P2EPePZ/sEQONDzAdPQcYnbdHfBj2qcPgET4cpwOFDGmsAflT08I3HO350BwUMrFMpcRG6ATqiE4CbAUHTpJQkNWmz2Zyfn11cXGw26/Ozs4vL8xeXL842Z4gIRIDYdf1ut7+7u7+5ubm7v+8O/Xa32263d3f3uRQArG5jiEmnxCyahzJ0wAFFrc5ISQqES5JcTUupF+PkgDabrtex94RwdDZDvcpodnkcbcMOEdpzfCfycwBmp6fmPVM8rI529Q+d1fmxHgxZxBC5ezW3Yx0xt3is24xDm0XVQbex9uPx58lR52bs6e24a8lRAARQRuMzAwpOV0n03YmYiRCRa9QRECITIiAhxAIcrhH8ZqqM1CRpmoTm6E7gbuamhACmZiqERIDubgpmjJSSNG2TUhJhJkrMSYRFmlWb2oYEAR3R2rNzSu3X795d3e/3Wfdqw67Dts3Cf/gvlnqDixYtWrRo0bdUSwTHokWLFi1a9C0VAsC//Ozv/85/Ai6OTdGOuDUnMLt8+aoVbVunKPfEjXCTUuMGal7UiAixBmi4g43UIuKG+64rZuAe3tu+74nYzLuhzzkXNWLpc+66noiJCIl2u10eBqrWWu+6zh2IEhpp8WHoEZ2ZVusVIKlBsSxAzapV4NeO3311/m53+Ppu+9k3d+92w92gB/XBfVrEflz0fsJtcPTQ1uxTdzctpqWUklIjwtWgi5SEAdgjeXkMr5hrZnMGCAex2ZR9gXPD8oOBmFWom4Vg+AixMODsY/I3eZ/dfPz1Uf5D7IooyH+FiA+LksFwhE3V20jSMKeTZgWQdjQCcy3DoDkDUZ9LKYpEKUkuJeh8PSlieQAAIABJREFUm2TVrtbrNQk3bbtm3mw2KaVSSsxJdPvD/f393e3tdrvt+97NYLqOoOYheI0KqbDsZNhGq6hPvfy4ntjooTv0sSfawSKke74ZyYOwk7HV3zI91SI/TdKoqQ/PAejv7eN7DLBwRLCPt3u0I4/RHM+kIzoRMFNiJqLUpIvLs83ZZrNZv3nz6pNPPvn0009fvHixXq+JuO/77XZ3dXV1e3d/e7e9ubm7u93e32/33aHrh5xVS7YajyMoPJbrQyRCAmJ0i5hhAkRAQWJiZpHIA0/SqKrX+ygmROy48iCmggAg+HNA3XF2IwD0vNez5AwvqvHkpDFc54El3SNwB2uRQ58f9PFIxHzJMSH7YRE/ACRiU1Wzul9m02KmdHwKxsOgqKurgjtQjQaq18CxxODYpyNCh7ieoi8MKIgtoDgwIEOtdMtINC1gAA/cjIQxHlSXcjiYm6tG8LcZorerlZsNXY8Iwty2DRlgJGibgRkhEDihgbAgMRITE/Gqadbrdr1ZrdtV26aUpBVphCUlEgHiYqUbun3uy6G/v757t+t7K4c+s55LgtJ3f/h/f/74hC9atGjRokWLviVaHNCLFi1atGjRt11//7/6G5KbdfdJvvwZrDCBnK3S2apFymJDYmo4CSUiTtISsYGRCLOYGiIRM43ZEcwMCCUXRCQmDP+ZGUDUEQMzcwBkUbNczAHUPKCku0fVu1g7H95qMARzLWamDgYIxSzCoINyHLp8GEpXbADYFvvm7vDZ2+s/++rqZ293t10uAAoQvs2Rs+EjioZjXmolR0gITITIxNykpmmb1AhL1M1TtSdR3RTNDHVhu+dSTLXWAZzRokDYkRLg7szsUEv5BV1i5si5MHdTK6pFtZjSuK85yx4Z1+SUHm3B9VhmphTMDCBo1+MUjhP27dWvjZMxcmwZArCMINs0YjfC3ekORNg0TfhCCbFJzaptpwNdXFysVit3H8uAkavlUvIwRFSLasl5OBwO+8Oh67rpdFRQOOZcI9IDj+0zue/o853bRxEm5/VkKyeqoSgAMZxmenqQxyEW31YADTCbZRl/e2wYP7lkHu9g6upEMx90nx75YWdG9vkHU+R2TPlUL/4xRzm8z4gkIm2TXlyev3714s2b1xeXl5eXF69evVytW0lJhBxcVbtDt9vv77fb29v725vbq+vrvs+qfjj0/ZCHoQCiY9iH611LRMw03moeUTZNagA8qnrWrnrNVcYxncfNA9oCAGLks0fFwNr4AMNjVb+TCI1pYcTkR4+ZsDlN5vFB8eBacohrdLZo49FozYn1NF3jT4117K029QiQx9MxTmiZFbfi5nAs/OgwG6vZ7qZWTQ3zWjaQSBATUossjgzACBT2cZuCpGvfZstKHN0cIB7D01WH4IAuJDWIo3qlgZEYIxuahIiJElMSWrVN26QmJUYUorZJ4aB3U0Rn8qg+qKUUtWxWEHm9BuZ9GTqFDnS/h//o//rjP/vN795fvP7xH/0RLFq0aNGiRYu+xVoA9KJFixYtWvSXQH/wox9pe+epBz4AkhMQQUuwWq0YVEzFgJDapmVJDs5JWMQMoqxTeNcIIezMML7AGkpBZgaOwBG5iUjsQOagFuvaFUe7oJtbXQsOEDwqao+hA7iBF9VSVM0AgBy3u3035GKQAXr1uy5/fXP/xbvbn32z++p6+/Z+e9/roVgGCBg9C3Y4krKRP46oDgHIwYGQOEmTmiY1JEwsQBy2Y61L7+e+3IpQCCnw0lRxccaVAEYAzczBWIlGz2F8P+yQREQUpQ7NrJjpjGUH8fcKhZGZcDzosWfulfi7E9XAVbWwW57YdytY8krTYv/uYGojJ4vScEDhVKwwd2J4EOkfQW9xpEVMHH0Mtr7ZbNq2rb5IotVqlZIQcXyZagKwlTwMw9D3/TBk1WJmQ4SvqBYtEedySlTH6moRmzC3mo6keTwfcCR1k9V0sooeySraiL1pClT56C00Bfh+WM/70/iZf0A/D3g/TguZQ8lHCSRPv46b5Dj1Mrt70B2nlAn3o+X2AaIHr4Z+Qoi7Oh4SwX8jGKFJqW2b1WazWW826/X52dnlxdnFxeV6vWraJokYeNFyOBx2+932/v7u/m57v93u9/vdYbc/HA4HMwfgfihF1Q2IGTmq1h3zZBAB6xSOuQMCsjBUYgvBxus8UyXJWKfQ3BEDO+vkVa6rFOpDq4JfxLr9w/P+YPGBH93oU4BPPXNu49VoEI2L0AxiD1I/G0SfZlfqcaYRsmOudL2Ysd4aY160uyOMqydizxblQsfQ7YhDAXhU2PAEQGNN3XAEYABBEho9yAjkY7hzLSpZ4uarJ3csQRmNCSCOCIzIjExIzEH8E5FgzIIRIyJCYk5JErMwCzMhCnMSbuOSIgJwQkzCAGBu/dCpZnTVPGjOakYs0jTQrgvRfd+Z8OBedt3ZoOv7/je+uvr9h91etGjRokWLFn3rtADoRYsWLVq06C+N/vF//Z9i3vD+k/zJv0UTVScwNmiJWLO4p6YRZiAMGqvmRCQsAIbgHOY6wrRqHdHdmYSZRaQmURCJCDMDRLAy6YhRmBmJSg2MhtVqFWkeWiw2YUEkLKpmVrT0Q0bERprdfj+UQixdPxz6oc+anbLR7Xb46Rdv/58//ulnV4e3+9w5dADDvLcT+Zi9BYFiwpdXoSoQEREDIUpD0hCzmedSghLPAzTiZxKZAjrm3Hncpm6moxnSTN3NwYWZmBlpyIOqBYMmJiEGALOAXzD6MiOB1h0giUQzDBwQefRHmxkShbNynndMT5HLoIfRKRHOpQw5IyIxR7Q3ArCIWSzftwDlETOiqiJCiObORBT1zQKda9GipkWEmZiIhqHPOW82m9Vq1TSNiDQprdrVer1ar9tV20R3DofDMAyllLu77Xa73e/3293u0B0CclYrKSJEHAqiqTKzSILqLcUxUMRjmMwi4sNimT8zO1YcV8/ANCIzXyoCGD4KNX7i9D0yhz651TP+NMZTR/EHdvUcAO3vP+RDm268+cRF4qcu2SkOGCKbN7CsSDIrqmXOoMcdBLn2mKKJJ4ZjSY00TdM27YsXLy4vLy8uLl6+fPnq1avI1thsNmCgRYch93232+2urq5ubm9v7+6urq7u7u52+13f9aXa8JnGGwYAD30uqrMGEBESkrmpmqq2bUtEHvNdZmpWsfE4r6NFAUCS1KfQOAtBRGBquUcSIHI3Zo7w+pg3KqUAADPX0PjTwTip4ljR8PjOFFSCBICuhYiRyUxrJI87InFKpnoaCzPW83uwugMB3MCskmFEQH484gBQl07Up1N8ZZpTmXPtD11xBCBAkfKcABNRImZkAChaom1Y70xAsLjO4yHKCASEgG6OAEzgrkHDV21qGkmpIQAGXxE3TIk5xUIKxlXbrNomSeJa9NXr4hVENx/GBRaI0A/D/nDY9/tcBjcld0aQpn35+s16c2bgd3nYuhuhHW6RW1f48R999oEuL1q0aNGiRYu+PVoA9KJFixYtWvSXSX/wox/p5tpSX9oeD+AIJdsKaCVCquAFXdGVEhPzGG5KEknO7qrFwEmkOhuRg2jRmK0RCErVhVPiVMIDDMBMSGQAqsXURKRu74AIhKSmploJIni8dvOixQwASc3MzR2LY1HsC97shm/u9p/fHL66764P/dv7/e2+zwBardAVOJ/WQ6tewOp4nNIWgtoQxz9IjCxTsEYcGaov2NEUEJGkGnD9JDA1fnWPNGYEcDBzwrBkVuI5q4BX/cbmYGO0a83QqIZBgNHR7O5Mk/eyhg+M0bKzaITHRsaotVgX7xMiMRU1NU0pjZkDo6NyDOSAGaz0MT4lnOk4MVwHDNsjjl2zCtaZubqhmQMQC1MSbttWAnmDE7GIuJqZgcNQci4ZAIZ+OBwOXdfnnM2t7/s8DG61cFycEED2uWH35G/S0ZMOWuNsx8kDGAvMzTo4lZz7oD6E5k6O/T4gPA6Kw1if7bHf9MEe/FlE+7EDGmY+20CCVp25oyu27h29JmkcL7bxu5ObGDAixYnIrLgpYLBxr0AXITVN2zRt27Zt07ars7OzzWZ1tmk3Z+v1er1erVbrVdO0XMNZ2AFyzodD3+0Pu93+/n53f3+/3d5vt9tctKh2XT8MfR4GNQNETk2N9KjrJkAfBF0H1UWCOncCq80GiYbuELb/OJNj390RPTKAUnJV13hwIUAtX+imQAxI4IrEWCk8IKKpAQASjs2ZjaL7SUnAKQVjvMfibWJCRDcbfeU2y4RHYvY69TQH0AAATHVpwzQ5YXVpxbRaAxGRYx7L3TSemT49VmsLx9N4ell/CEATIAMIQEJKSOw+Jj6jAxRXn561Y2cQgME5nMtECEBAzBzZ0CLEhETQiKQkIkLgArBJTcskUenRzbQwkzAyY0zrFVVwIOScs6mhQzE1tzpDweRUI6pF5GxzfnFxocW2w2Gr2oN2ORshaIHh8OM/+uZ9/V20aNGiRYsWfdu0AOhFixYtWrToL5/+h//2r/Nu0+y+sz3/qauRYwMsYKumIVfUDhlJmIndXU2blJgIwXPORYs5xP/VB2B3V9WUEgCoqpqpW8mWOKXUlFIRSJhYHWpsRQW7gSqImGnoh6h5GFhWzUrJJRcWQaSsFoiJENWgqBukAtwbf3Pfv911V/v+m5vt29v9bZcPakMEQ+NIao4MupKbWKaOPi3Krz8dEIiJEzctczigadom/JSgGRycBMaoivG8jvgYYFa+DCIUwKfs2NgSoaZqALoZVAANdQ9I1cHtlXrXFnCkNlsAaKTR8Ih1rf2sHSei0Tx4ZMrgNnqrfcTxRyPo1KWxYFiUKLNjti7UeJBYRz9mfsTFkFJSq+LRv4wARJhSEzRcJDVN07ZNIhEREYZwchPmnLuuG4YczvrucMh5CLqtRXPJZm6OJRdVjdwDPw4wAk4obALQY6eR4GF5ySes8j+PHn73SWQ892EfQ4Tfh/uOtdueY4J+1PggkePVZDgD0LUJUM2q4ID+gL/jHOaP4B4RmMKwiyIkzCKcUiMpJZF1aBOoeX12fna2Wa9X7WrVpCYxs7lr0WEYcs7DMNzvdre3dzc3N4du2O8O9/dhgd8NuQASEY+XmSESMjEnr/Mi5u7oDo+qRAIyIuJ4H603Zw7Q7Xfz+3Bk6wiEQX2RGdzAfLqVoigfIgAxAAQmPrlmJm47zh7NPnJ/opho3XK6/8OtPX3RwcERA5CPk14j2p5d13WmJ1ZC1MvM3MzHcqZY/fAEiFZZrZl6TKCZjTf9FCYz9z4/eDE2fPwpgILIHgAaCRy9xm44gKEfW+keU5JMxADCNAPQKCyB0UU4CQkTITEhMZE7A6xEEhFDpNCrlozgjM6MYB7LMdwBiUvObs7IiACM0nBqmqZtpBESRqLV2UW7WlvR6932fhgOfdlht7+V1dqkgR//5E+eGKlFixYtWrRo0bdVC4BetGjRokWL/lLqD370o6G5yXwYVodmEGEXaF40/PrlBbsiODGLcCm56zpphJgAIOech6Hvh/DqAUAseGeqC7HVTM1LUSJmklI0NgBCdy/FxmXgYf6jYgoAwtwPQ8nZAVJKwtIP/TAMeRguLl4Qye5wCI48IghDEkdRkO1Q9tkzyPYwXN3v//SLm6tD3gH0AGXC0DBGmM7oIHqtMzbR3ZG+EBAjS9s2obZtU0qRTVGKRgxy0TAe4imx9SN/NoP/j73395Uty+77vuvHPqfq3ve6Z2yJhCRYqQM7IwzBoA0wcOLAIXNBMCYwwMCJY/4PhgMSkCXAggIOHMgCrHQSQxHhxBhABiUTBjVjTne/fj/urapz9l5rOVh7n6q69/WQIaf7fPv16/vq1vm1zz7V933Xd39W8j2Uzay2piIbmrZDWq+5y825jGETU/S445VrjIhELuOexZERRzNzj+QRvLjdYQldpQES8YSPxHCvrFY3Q0d4E4v042aa0vvmrBLmHp4Vhdwz3BDOPSUfIsLCNTtPumeUPtyZRJiJOdseatHsxSgkyiLKZZ6muZRJpim96fxzoQATifCyLM+n06ePn55Pz5fz5en5abksnvDoZtcbeafu6/UB/PwPr69fo78WTaNve2PYflf8GZtx2eOZ1yTydyjos17mdx76+ioJQDwO910uNgXy+YjYmjdunOGbigyCibToYT68efOQzvLj4+Pbxzdf/vjHb99+8ebNm3mep3maSnJ683OjLcuyrsvlcnk6nT9+/JA6nU7n8+V8vpxOp+fzWcoEcGve2mruxAxwBCWdOecbEW04m+irCOSWjZPquXuSHNh5niPi3BPQm40L7lUlatZyrwnWkKTKABn3lo6yhrlT1oq2JodEWYpiEZL7B+2+uyD654BdM9A9ld6j47E92v3jdODXc4K8um3mloWEm4x8DIJ+eHrW7tEM5rBk6fTPhA099MpufhV8puv3GZAkPmcgnIgRHMEIylaEABMXVorrcgkmHI7HoiIEYcpfSKpPoBSdShnlKPFMoEeQR2bTwz3cso0hIQShTHNRYSYQZV9JFVFNxvzhcDgc5+lQuDAJl6IkZAE5vvl0Ov/qw9MSdqp1+fjpP/n5X/y7/+i3vpq/+Fd/9mefeyZ27dq1a9euXX9ztRvQu3bt2rVr12+w/ugnvyPGCkzEHvRY5rcP849/9GUR5bB5LsoEeOaAA7AeQuxZ2VwmHhG1VjPzzkbocF73qNVaa80suRHmnkHd1loAxGTZQ484ED0wK8IsrbXsRXg4HgE+X9b08DwMABE1i+Ywp9WxGlbDaamfTus3T8uvPj7/f5+evvp4/nhpa3QbOlt8xY1nR7H5MsCdB0OZkxVRVRVmnbKFmqrqwA1Ha41FiOSmOdgtAxrerSsi7lwL2pbGJ/8UxKNr412QevhlSXzeksvMfL8wvx/RN77EeOXFewAgEbjJDXA3MxImkc3zttbCfVBBeIuXxmhOaOZAsMj1OvPQHghnCnQ7j9MmatYylzxgHcEs6bJtDf0ymSvcmdqiooVFIcIiPG3SaZ7KPM/pD2bbw4hozYBQ1dHVcM2bt65rdrHDjTVvySPI7PTnnoXbISO8sv9GdP7Vdn9tn3rskLbelq98v9s8vvd8/qvzuP1D3HnQfeZl3PYGsHDXv47QDcwOeiERZhYmUtVSyjRNh8PhcDiMWS+HeZ6nqczT4TAf5rlogjREbzrDAaitmXmt7XI5Pz09PT09nc+ny7Ks1S7L5XK+nM6nuiZjI1pra2vMQiwRlM81a4lAWICplDId5ltTGOjdOQf5Y1tOcMO3iATm+GE+CHOWxNz8mtxnMIuqWLOtJyfRFaSRHjBFYoUiic85pBHhARUBwt0gnatz1V2rQCCfEWt0w+EAOouchfNUqTNhSERA+bmRTz1eaHv84zY/3UHoEeH5QYPackWFJ07kLu986z5/Z/AZAHXoc7rPJCABE0EApmCQMAkxMymxculUGfRelEWVk6+O4AgKZwIDHMjWlGlAC5Obw50A6X1Zvcfts+0tIIQiPE+liAgxIVPyMhWdi85J8CjiHGlaP7x51MPDpdZ3z88fzu3U1vXcPnzyH9enx0+ffuurj3/4+mp37dq1a9euXX/jtRvQu3bt2rVr12+8/vl/+w+AUDbio5b5xw8Pb968nacyKx8nnosQAoTgjihVVUS4pRtCRHS+nFtrIBJVEWGImddma9rPZpvJki7KsiwenqiNTO4lMjiXVwOcFmd6De5YW+srzMMSMLzU1po3Cw+qhktt56We17YG/erDp//3V+/+4quPv/pwfn+p52aLhREc8HT5rhG/z3i1PX1MV2svrzlducM8A5RBbGElYu+mHnUzHkFpQN8hOIYxHJHetIcTwCzCDKZwmHniLrZT8vBkZ0R2JxP2YQdTZh49oSB5ssRpUvcGa4HhXG/+V6JsswBAwiwi+f5RSaCbZoY0+NfJcXaziOgw6YFSGecDIbLWwkNU8lo7upulNfNwjBNEpwWQNWutWm0iAmL3IAqiABnCA8FCKlrKdJwPh8N8OBzSED0cDvM0lVJEZZqm4+FYa12Wy/PpJCKllOVy+fTp6f379yxZ7aittexUZs1as/DeWnEQcuOGLLLdys3THxHhnp/euAufDxajf+v+h+Sr6d1ZCp/bCjyyyNGdvLgamnTzn6sXfp/UHgYobTzgbDqZll+ySRjcX8vkr0zzpKrCMh/mw+H48PDw9u3bt2/eHI7HeZ5K0eN8KKrElAZga21d61rrutZ1WZd1QaDW+nR6XtZ6OS8fPrz/9PHT09Ony7K0Zr0FnkfrdAtmkRiVCSJmUSCIk8gc3pyV58Ph4fEhawbu3j3gLfU8mkt2rsUoiJibNXOzwzyrCgCzyC6avXCRVGLVm1oOAbDw6EDzjgciJkTUfs651gHuoaIguFXceOBj+F8qIsyNxmOYHwfeLBAi4u5uzsIAhePegObr6fU7jdtPqxhXnQY0PCnPAXNYexWe/8ypfcaAHjCajssASiR8I1eFcHeNCUIJYSIhFmZhHcgXp20mh3sY3Cmc3DXT0JF1J2MiIRKBmxNChVWLqgaFqs5TyeIfIYpwUZ5UVUVZ8h4xy1RknnQuhRAetrrXcBN5ePOmur97/vRU/dzqaeX29/8v/Pu/u3zz9n/7N//m1Tjs2rVr165du34ztBvQu3bt2rVr1/dBf/KT3+EoxWSZiXkqeng8TBNzoVbCVCBCVFhURQVwERFRYRnc40wXMjOJiEoJh3m21ovwYBFmTmfZ3RP3HOljmnVjJQCCW/YyZBGWRHM0g19Djx5hkYFJZtblXNdqBj4t6+myLmbPl/XptHy62C/fffy3v/jLX3zz/M3TcgFWwLKfF90xeD8XGd7c5+uSeWZmUVEVzp6MnLlm8xwNrrW5WziEBUTuEeFEHYgRwz7KPQFwNxUVFSdYbbXaSPghU83pJo/IY4cb94HoFOvIP2ZENNOsBDRzJiImdydiFRmH3hAcvfljvrJRua/XP9oh+mh42MkF3L1TG5Ztng335mwhLJHJ5ogcr8hDhFO6oB3y0a32jNQTIKIRZt7MGiGI2d0JUNGiKsLpXBEwH+YcGWHRooepJIJ8WZfHxzc/+vLLuUxEMG9v3jxokVZXMwMwTZOZXS7L5XR++vT0/sP7da2pta7rWpu1GG5ea9ZaS/JwXisIHQhOFN17fyUemA3hfl/iNhRL29zbYuB5U9GLCFsZw/oc3ILMPU1PMVgj6SZTIO7i82AmUVbRTDQfj8eHh8PD40GERaVkKeV4mOdDUS2iPeesUrSUUrSUqUyqxfsqB1/Ol+WyXC5LIC7L8pdff/30fLqsawQul8vT01OWT6o1d3ezVqu16s24lCwtRI/idoKGqlp4bS1LFDLl+gLJtQXuIcIiKqp9+K0bzDfCoKP3nSM8Ge0R7u48zOEx30cxYSSogTt/t5PW897l8zE+HMY96usliCWD1q8Z3vcZ+e0LvxYk8jXf7l/ytfNxvmtUeDNhmHqLT0pURS+iUUSOC3BDdnZ4XKfWX6EbD5r6GTGghAJWkII0KL8QFmEhIlEWpjxQRrkRoOAxUb1zqJkjzKwqixIXJiVIdnDtVBhXleOhmDWiOM5Trn0pUylFi6qWIsJEkWwXIgiBOatYRAFlYooIW5ZlrQ0s0xc/hpanej47qvnl0lzqOl1qOfuXv/rpT/8aQ7Jr165du3bt+puq3YDetWvXrl27vif6F//od8/EZ5P5sTKKOAnoeJjnouJV0EiQoTRiT+CqqKYv2T022sQZmSaWnicdYcy018wsvY+MUadp1A1oD7ere1JbdfMBxA0CgmCABTzgQFtaswjitbVLbbW1ZbV1saXh3fPlF99++OW75199PL07XT6tdraBQSU4KDqGdTva9hV99oecTkfmRBcLq4CQ0e9OdE2DiNJfTuwHNussU8lMI4+avc5AgXRe/WpAD8Mzz2okQLfudXRzSj0Nnf/wuIz0eN0th/315Wyh3rjN6770v7DZd8wdvHtzhtFTzURCbO6IEJF+N3OhPKsTIsLdmCVz7p3zMSKltKV6KRBZnPAEXqfVJmnmmpu3CJ+nObPzGeyVBPgSRfjxeHx8fDOlZS308OYwTepuzKSi8zwzS1Ia1mU9n0+jU2LnNFjLrKwluzy8J2pr0iXMWTg8evkkIi3mfF9CHmxUAjLWatZ6xrqjQ0JFiXnzUzGSvWPq9ZwvM7SoCJtb3p5MnDIzxbYQQUQE6dGXiQARKVORnnlOdjEdj8fDYT4eZ1UpRTM5LlkQ6uTgPCK1Zq3Wy7JmPHpd6rIsl2U5n86X87IuaxDW2t59+HBe1mZOzLXW8+kZJHnzkDPDnYmEWbTkEEU4QMKaHm+WE9y8e+pCaW4G+mgxDbi5Nc9o8uY2d8e5G54RuVF3YId/7/cO7A2s49UM73T4kSSn24+Bu3clNDtIsjmh4TaRfX1gBpRjOyZv2fmXD9ZYnIDbD5x+oGuRIW9jB4WMjxIPd7c2KEjen+N7rNBnRuDVOWw2enY4VKJCNJFMxIVYnGSgi3I3CXSOsJzVkatFfLvqTo7pCyXgkxZlFkIhKgRyp0hyjkyTHuciQqpchEVEi07zzEyByMtmDmYhwL2FO8JzvYUy5woQc5MylekYPK0ez94qqMKs2rff4vgQOvv//H/sweddu3bt2rXrN167Ab1r165du3Z9f/RP/uHvSTFmigimbPdEhfh4nJRAvnI4U3DpGd2OSdbibtExCxQgcwOYSUUKBt85YmSB00LK7OGIMm5J2/BwCzNLbEJaPOHw5mEGgIQhvJqvtS3L2jG4BAcM0ZrV1drqq2F1ukC+PS9ff3z+91+9+/qpvr/44lEBC1i2YANu3J8tEvhZAzqSYirCxMLMh4ejllJbNfcIFNWN3JrmTMaFzXvKG+j550CkQ9fMrBk6dba3AOwH8zDzNKttZEVfJbWvp4th2AEgFvQsrfUMJ73OJPKwAAAgAElEQVT0oBM7ndxniCJLAiIvLzyzoh0PzQBYOOPJebvT7lTizESrSniYB/fAOhm6PZvo4I3iCyACZlFUQVjWNa1kb83ckgZOvXthxqXdzCJ8mqa0NdOyDDerNTxK0QzaRwQzlaKlsBYW4amUqUzTNB0Ph4eHh8PxoZSJhYvKhjNWlYhora21tloRUNXW2trquqzrutbaVNXMzqdzRHSQiFsz62jj1mptAUjRfIjWdc0Z3lprrbZm8zyr6DVVPczfbkkjcm2Bqh4f5mnSas0jiChPU0RykUH2aCylIOJ4OL59+5aIpml6fHzMVpDNWq21tVZKya1UOTPRtdWkZl/Oy/myrOvSzAh4enr6+OHDN9+8CxATXy6X59Pp+flU12bNI4JEgriZBxGYRSTCrTXWwiwj2A5zV5FSCoMQYd7JG6olnwsauJgs25hndz03jGaDEW7WmkVdwx2iPTO+PaRJ6Am67a03GjveO7DbzB9m7ssne9BK0hB+2dxwe1PPrMcVlMGv7eyXvSuJiJXwsifo9u7tee8bXh//2Az2SCI7b1Wu7LlpzZq51XDrxa0eg79la9wc6sXjP4z2bSkIExWmQlyIJ9aJpZCIg7wvWjFvMRoPAh7jQARWaH725+gyBQAVmUqZVLMD4Sw8CWX9h+DHh+M8lSL8+HiYi5pZKVLmqZRi4eu6WmsRTpx9blvG6s0qIYryPBXrWHr90Y//1vH4+OHp/GS+gJq1YAuTtuJywU9//vPPj/6uXbt27dq16zdKuwG9a9euXbt2fd/0v/zkvxQNna1eBI2M0JzYY2Jib2hnkUBYWjAiqqIRHdY6TZOW4hEqk8q0rNUjhKVZszRhR7ovTcjWqttIQUeAyFtrtaW9qFpaM3cPgEFMxAGPaGl4J5jV8+BGzGCOCDe4wSHNeXUsFqdqn87L10/nrz+dvnlePi72VHEJVAADmdCXwH8e7JsKwmYEUfScqQRxMg0y35xmHwZGo2c3B8wiE59uDmAqpVkzc1Ul6tnwHEbcpKYBbFbdGMCrcuiE06SijJD2OOqgD3Rz/yVlpEcqM5oeaSjzS6vsjtGRQd1MNnoPmSaUo4d/A4n7GMnirfnbdkDGLT+533MCkYdTd7sjvCGMRAHArQfMweEN7qwFhAhn5tzCWwtzyu5yInktzBzRCEEZrhQhorR3D4djKVNPsauoylS0TGWeJtWSGGsRmaYp3cZWmzBng760lTOOLCx5n7O3YfZfY2ZVTc7MWhcVLUV9FFSmMqlqZoez9qCqpWggywGecVcRmYpqURJO+nCEm7m75S1Ll1pEzIxF0mVO+9LN17U+n57Pp/OyLlOZW7Pn51OPpQs3s3Vdnp9Pp/Plcllqre4OprZ2FEn6tT0EnlHvbpQLmAdTZRjod0ne7pumqy4sFHC3tTV3V9Exq4OJC4sNzEcMoMzG3nbzVmu0SgDp1AEVPCAWvh08DeTgrUMhcPs3FNpc5Rvwzgvf+Bo27u9mefUgYJBkRASgrVXgy/282nOEffenyrbI4cYgppHsBjaod74sRHCvrdW1Wq1utae/r3yRz7rPGAb09eS4L6gIQmRmWYiKMAMcRID0xoM9AQ30e8sIHhuCwDmgHkxgQoKhmaAqRXVSLaqlaFEpRELEiKnIYSpaihAhnLJHrIeoQPhSF3PzXBVizazlreOe0QZRiKAUKYfD4eGtzsfn8/q8tiQstUouFUGg2IPPu3bt2rVr1/dJuwG9a9euXbt2fQ/1J//9f26NrNKyorCtwa0RPA5CAqd2DlvhrcORs6tY+LIsh8NhmmdiJggga20RYObeSywjzMCAdXBrq/lYzZ1g4oxEWiNiVR1dCUko7V64e3N3UBDAyJRlmCUuNQLucIMHm1OzCFYHreYfL+u35+Wrp8u7c31/8feX9Wmp56VZt4hoI1HcWKQvdLNMv2cImVgOx8PhcHT3tAJLKcwcHhkcFeXNVEoDutZGwDSVNGpVlYl7c0IPD2diUOcsg2jzFuMV3TWtwL5Cn8bpD1oBM0eaxUk4udVNfpNuktQvQtYBJGFi+PP9u+mGwjsrI9G7QGRM2wdzIq32buyBqZvxaUL2Vfbd1O4R0xxdp/AgBoHyEETEArdwh0h6ZxsSG+GJQk6nOWnURBRmgUCnUXTcCgGlTCxCBE2QxUgHz/M8z1OZpvQsReRwOJairbWplMM8TfNERNkuUli0M9AJA9It2hcFWLNmzd1K0UnLxk5gYha+Db8nVxzbsADjyjJbrhn0NrNaW63VRpo+CeyXdbFsFMlibsvlUqvVWi+Xy+VyWWudp7lVe3o6m7l5r3CY+bImATtpI0EEN48RBu6zgQZ5enBT0OExsVUgtsLNtW/jmEw8cC3LuppZz/CC3LMHHeeEv/qnA4ENJg+YGVqWEHS711loGT4r9zUD3aMc7xlGtOccG+RuIvIb3szNM3Ql0qA33HsZGQ7O0oizCHXi+WcQHPFq3x72qvjzSnF/uNuHMLYwNBiB5MS05q2F2xW7kaWu8fsr0c0vELpfzwiOYAQFmEh5LEwAKEABJWKAQQTKag8ni5kiPz8ExARGR3Mk20WYpqJFkyLDKjxNSgEOCGEqWopmyt2tWau5yoGYHXi+PFvERtVBuCa7XLgn+RllkukwPXz5Iyc+nZf3l/XSYq1e3Y/2xnVxrbv7vGvXrl27dn3PtBvQu3bt2rVr1/dW//gf/S6TRzB5CWpGTGYaXtjJFwmjSC/LHh4fI+Ljxw/TNB8OB5WyrO18qaXMxNzMVJWZw2z4Q8TCIuLJEr36WTSVUlTXNdHOwVJEVVQz2yfD4HEm87auy2GeVcSaRVi4N4uay7VbmCEMohOLVDNjXVner+39pX57rr/86ttffv3+F19/SijHwHFcM4TfZRqNN/SegNhcOyIWlVIeHh6LFg+/LJdq7TD3pnm5ORHVWgOYpukWBBxBA2PCqkpMa60b/jWZ258/n4jeyHFATjAsrOzO5xH0KgGdacl0Ez1BHICN/WxvMzN3b2bbKx2z0Mxb9dbyYADgDgRYeg+0PBN3MIOZtDAxg/3mdjOzlpKHY+bsXUjcUSTu2WlScnxUJEnNma5lhnvfUIWZOX1hTjwIkTBn5jI6ACaD4P3q8qKmqahwtrAjwoB7S2vVWrXa3r59ezgeW2vdrU5HjTNknYe4ep5EJKXjPMwDgKpsPSszs9xadQ8aFGxcfedgxlYwcEuHP7borrs387p2lEfSvd390/PzWmtEEFBr/fTpU2vNw0VK3vFSJiY2oyAy93VdARKRUia6mS0RMDcARXW70+bRzPKO+wBXJ3GYkUj3sPFQx7XfX8ba4SOK3mqz1sIaq7KqNcuU+nicRg89HxwJVTCDGGZwSzgPiPuLDBEhliRjp1WZYfsxrh03b3ZtzkjjKl4/1yPQPb7psTnc28PSs/sekA1B8VfZyrnvNMw/Q/S5PQThpo3kq4T2GByrCOsb9yB3H7EeSf4O0TX+TAAxnImYWAMMCIJipKH7OxgABdKe5uE+E6DMwiQDBs2MSeU4zcqdjq/CwlKES5FS1JshnIWjNXKfS4kE3SyXVpdmK6IXexAw90tbQSRFjvN8mKfDPJVJi4qKFmEVJubD48PD28elru+fTu/O6xp2aWs5nRq/jZhKTH/8p3/617g1u3bt2rVr167fJO0G9K5du3bt2vU91z/5h7/XxNeZp/UsoUr044fpR2+OXM/WFiaUMpGIeSzLRYRUlLm4c3MOJJWCc8V6KdLho0SZxVTVtBrXurq7Shnk3+imIZiIWYXAGE0DI4KEPbxZ7dxfEssWcp7RUbmc19YMYCJxoDWriNXxYVmfVjs1e//x/O2ny7efLt98On376fn90/PzWi/mgw1N3WW+Emdv89GEDEVupk/ayMzEojqJKotENiZ0E2ZR9QEOsB6f5M2A3ogUaTjmsNS6biZxBlGvP3ptdjZz55DksGzp03BEsCqQvvav+5ktkqccEdbA0sPIA0HbDcXe266je63naS1HRkZjQRbpuAYRAsI9N/Jx1gmRyFw8b8naPqTDwXT3CBEmkLvzaPsY4ebOoyVbs5ak5rEFtqQzOlKBY4t3x9WHMxtkkEj33jDCvsM5NWvmzebDXLQ0a4hgJlHJ/TMzEXwQzMMjXUotEwtjUGZUEwuRDioxcU/aMhOup9pvZZ58j7mHVTNLzEiatD1uHFe5e6RTbe5hPrx1cw8iRgznlphIgsgDaeu/ZCH39LIj4QxMoHSD3Vvbwu99trPAgyKIJQjhcU3e33f/22L1PSAf6JwcvwkiMxFz9pnEmHR9ciRIOz3ugWmOK2aZEDROzXLtQE86b3az39Rd+knaRqe5jjtoLGiIxFATX5/NnBWxcWyunwK3RZ3Xwerb/QN8t4AgFwJcZ+R2SUSUxaqNVpRrOtL3D0+q+/0BNkbHeP3qX6ezfP3FSFhP5EeJBBggZMwZzETR2RoZeWZ4gjg0H3skW4M3fAcTFeFJdXT+5Fz+kPcTBGvNzQguRIXl8XCIiNZqa2uEEUXeemut42tKKUV10qnoPE/zPE2TinBkap6ZZAotn86nc60rYTV7rvZcPx2DD7X98Z/+4vN3YdeuXbt27dr1G67dgN61a9euXbu+//qf/rvfk3Yh1DkOs8qPjoe//eXDm4eDrychzPNs7uYR8BFmFOaZZK7NACoqtVYgpqkQUxA5opmZtVImZorwZV3MrMiUXs+Ai0Y2e2NhgCMQ7mZmZiISBA+j7GnGas1ah+pORcvz82ldW1qQ7lFbW81Wa58uy2JhoNPFTpf2vPo3H56/ev/0l+/ev3s+f1zWS7PFowY29qkDAfDw06i70nDOqORtZJr6OnURKUWLEqPVJiKllI7UQDeKt6hxz18OOAlACYiw1tJB7HHRdHRiA2YAaWV2x2oDdHQbMiIoQ9O5E7ywwCK8G6kdEGIeZiTKKtist86DYFaRhEdw+sK2UYCZWFTS57w60clHdk9OxYaEzkGg3swxLzava1C4PVprZjbPExG1Zszcc8fh7p6h8IiotQIopSSYojOAx8VFIHpLyC2gntgBJFg8ba8kUOCevhIe4eFmIpLM7qAggghHhLX+uoX36Kx5hANRppmIM0pMRCLZJvEKrCDmF+dJBHyuS527u8VGeUjXW1Q7YbwzoUOKJi/XW2Pm+XC4Znkj0+0jYI6r5xyBsKtZHH1iDJgDEzG5R5iF2+by9tStlKwkXGsVNBzVGBHmLeB9nal3FZRBi7g2WOwO58B6jFIHIqKZcYznjhADQb5NaQ8L97DbFPG4TtxSoQPYsBXjLSBkoj496Ax0q4R7dDOaQATbQB24fQC34cMY3vGfcfkxlkrkW7fnb1QUtmHalkj0axmJfXRbf/v91WXeixKzgdgMaAYEIJASjzhz0p+RVG3OSh0RZ2J7MLUFpERCVESVqQ9V7/kaQDCgzFOCZ0SJyBLcvM0+T1aPHabpOM+HUhBuZhlnF6H8n0KrlZhL0cN8KEVYiJlUpUxlnouomDUQqZQW/O3Hp/drc7jB2sr/+F///L/4j3/77/wH5af/+i9+/cjs2rVr165du35ztRvQu3bt2rVr1w9Cf/ST3zmsXxyf/xZ++y9V9IuH+be+fHz78CAU8JbGFDMjzK3VxUXmMj00RyIc0oZwd1FhlWbtSpAlMHNt1TrngRDUO88xqRQRTa6CmdXW6rrWWjuaginM3DyJuu7BJPn+T5+elqWmt+gRtXl1q9bO6xLEUqbzuV5WX5wM08Xomw/P3zw9v3t+/vrD08fLerKwkYP2q+FEuDpJcPJu8MQLS4pBlO3jRGU+HEWEibqnS+nb5O4oEdYeYe5XBOtI8maW0zcDOg3vG7e6e9abN5auz6BOiFzhwi9ik17NzcpUVLXTLVpb11qy911nfgiP+OdgGxALE6iZjcBsTyT3o4/TS4SEh6sIcDWgfZxKd2JBiQ3p3AYCgbLGME0JXDZzR0RGyN0t+drmXmtFQItarTm1cGPmud8Bs3O2ZMzWB0Y5rCFAWsLR2zASsfAG68jL93AWZiEQhbm11vfGjO4vZ/wcZSrElP0YBwgiWxSOrnk9CTtO87sxDixKxNay6yDSg8+JgcSFt+bmUhQgdw8zYtJ5pp7kHWZ6DzLb3d4JtHX0u57JMKDzyfK+A0roRJ9ERNyrGiwSgXADMcU2zwIRoqKqfHOlvSaRVz+a5dV8aK8TmTZ8c55DHggRFPzy7x3UfWoCgcLNfIBiXljfSIOfKQgvHlT0agNk8G02bMi2XgHjlH7NzbqWT3qEvDf5+67qAiKRJgAwqiRoOe9bX1uAjbLdnfYNfuJ4/ZHzYu/ji3SfC7FSJprzs4myvpfkjZ5rR0ha1cRClJyNUkphEaLkLwPe6lrr6q0xQUUQrsxzKVt6PQDAIxwUvW8lEYPePj4+zHOrNUsab948alGQz/NUijJRKSqaH0S11bVZAzkLz4fDNE8sYiS12cfLUoNreF3t4cv6579c/uLry//5F19952Ds2rVr165du74X2g3oXbt27dq164eiP/n938fjE82Np/o4SzlMD/P0eHg4zDOFk1emADzMvDqCiTScPGDh6IvJI+OEHt7MWvqAw2z1CPfwbmxuuU+KGDiOBA601hI9DCDTdImDAAAKj7R/lrW2lowEBGAW5tbCDRlvRWtohuZkXKrz06U+r/VpXT+clven9dvT8umynmq7eLehA4ixVL8fe6yTzzPtX2T8kIZDzFxKYUozWllV8pVEGzNv4VGPEGbcY2rT2c2scUcQfMZ2ekEZ6EiCQCgLxuYvtnFzuGsp6TK3lkWCSKougDSge8u7LSo7oBPDnutx3p4BvQGSWHebXUQIZO5b0PtmnDo6OTELffOcDO6qigxRu2cqfCSgiYhiEKuZOQ1lVrmmTjeSRU+gEghMPEAC6I5wmsKiDBr25JaZTmd/ZKiZSPql0fZK3r64epMinHZwXqFwj+1Hn4nDYx8ZXhHJi315Rzs3g2/vbT4IybmmzLibb2wHNyeCljLizGMebgSMF7rN3vYCxo0BPVgfiOh9/66zqI9hnry1luMAvxly6tPoCoO4DmX+EQF0cMa1B+DL4DSN3+nGxr3uJvscpltunnSRz/nPxJRdN4FXf3nJELuwJALEMnpMtL03L3ujq78YwtcvvnjSxuMxthhvuZaF3HN00n72Zj317HG3l4iA44b1/F0GNI2L5MF0npi1z6UYvQqReJqN0SEgAZSlsBQVZWZGL+k4GCAKILxVt5bDmaFpZZ5Vw6y3IRUWYVFINg9Mhr/IpKqs4U4EJtLko/OYO+5pW7ubeQ1r0zxpURYp06THN0b09Hy6uBnIHS41/79RDv4//qs/+46R2LVr165du3Z9f7Qb0Lt27dq1a9cPS//rH/xeKRHaJj+4qIo8HsphehAGRyNvCEPzaO61hz7BEj0RSpu7Wmu9rEuMRGwugXcLM3cLZs4F3LW2tba6rt2t5EQTpEeDnu10Dw8WIWKzBgzWQlCmKwPp54RTSJFmtqwVIRFkjhZUHauhRtTA4vTx3L76eP764/O70+VDjeph4dXDYmPFAriNRN7nEenmd3TPh4hknjNxPM9ztgfs3fS6iZmkEQp0pHNGL6n3f+ueaFqB26G6i7rlR0eS9HUC+sV9pMHBIKLwqLVGhAx+sZmlE13r6oPVEBGt2XCEsQVXbxPWadsSqPvN7ioCIhsG6I1HnBeFLBu01jI1Cep52/GF96ArS4aNkxksKtl4DhliBVjkRaSXsnLQEQjdFGUWZkJE21pigoRE0/3PPof97ZT+KHVAcQDBzEmdxuYm3/84fDWU84CBwViJEcImANYMESV7stkd2DfPucMwRHL35p6QcxERzThqB6kjwKDkfqhoHo2IBzY5U/y3BZK7iXAzk6/3iAijc+PdZEtrlLiPZc4cFu6Otfc9def6fljMbpHM40q3ObxND+oXn0zn65wem1zjxtFPVajH/u9m2HaFY1Ji3O7b7+aTslUmbKTjt1eSxLH9cezxZi8bogQAwa7dLiM644K2saaNV5LKdLx3TkuE49rw866KsBnQ+LUiYINs3BrQQhQBz+aJkfCNyH6fDFaCgJWosBTRSVWEGMj1JdFymnX7WwiqCWgPFZlEJiFvFu7M0CLTVA7HaZpUlcuUTWTFzNxCWbJmUOtKRFMprbXaaq11XZfWVmawQIS//PKL48Mjl8lJqsVzXWrQGmRYXKtGYaI//tn//etHY9euXbt27dr1vdFuQO/atWvXrl0/OP2L/+F3P/Df+XeH//Q/e/5Z0xJVzJ0pDmVSArXV1rN4KKiuFQHRqbbazHpilsm9x/2atdbqWqtqES0Au4WbXz0dgnu05hl05NG9MCJUZCpToC/aJqb0FtNiZJYItOZgJnCkJToi2ABZc2vemjeL6rE2P6/rua4uU6VpjfLhXN+flneny/un0/vn88fLspo7aDOBRqPC1I0HfWdAUzZtgzuJ5Np8UWVJyC2TMBEFaDPvmDk6l8O79eSObl7Ki5++wt3Nu6+ZYUJ0Zz4iWCSdLrq1z/K0RpI3bTBrBqJSNALu3lpjZmExa5sPGO6ttbT5WJV7zcC61dtllJFgEgBhNhohGpCerKSjZm4IRyI4iCN9XiHES0tXrgzocDciVtV0gWPARjrzJC+Nbr1BimtjPYoI80yaR2uNRTrSNu7sPjOLADObWYR3a5vCzIhIRDuK3J16HpiSUbxxRoBEkye6gwdeJjE1MGtMTDkIIBrDeDN/OiDhtrNceJiZqCQ+O6KvGsiZ1M9ZOLw3H6RheGcZKHrNAC9/gL9a0FsCOinbyVC5PoyZ0w8LHlhud2tLJZUtMn0TdX5hlkbcRHpvmDGAxwAcY3invm2UJQ68cJU3/HQMnkcvSd1XBG7rLsODxgslPmUgOCLBF0zEchOW95d2890AUj+Z21UA0cHr+czeflIkiSQh4+HW79eGJNrO3e06KftQvTag++3ctiIiZeFI2oZvDOicSAZPOMvWWlBZiqgyK5MEcUQCaBI8HWHkoED/5KIoKqpCCGFSFgaEqDALkzKpihaZ5vLF2zdaxKO55y93c2tmrV9UVrwG6sSJYNaA+OLt4+Pj4/HxUVR1Plazd8/Pq8Ek1ojVlsvf+7eH978t9fhPf/bnL2/Erl27du3atev7q92A3rVr165du36I+sM//MO/u/75m/r09sNS35zM0CycQGaFlb1iuXBY1AoPdKco3DtLt0cEOyvCzH2aJi0TSAiciNu0YzLDa8OA7R3YEIkvmMqEcEsDmtBb5BEAqBaAzALEEVRbM3OPYJHsbmbN3RxOS61rNQOWup7XtUJaaMV0Wv1U/dTqh6fLu6fTu6fTp/PleVlPtS3mFclsGJ7TyPW+HKmMbaehg9GLLBOkI5OLbIAW8IQ+Z2q2W4JdlPBlkswL083SdbNhLY54bQCRF8v00pIDbk2r4RWGW2IuOo45PWVQb5XGBCIOhJvlDWXRpG+ktSrCwwOMbMdHLGkPY0Mvd5N8+Hqx5W1730JsLOkXXjlARCJs5ubGxCIiN2jpEaLfMuA00rq47o4AIo9wc05YjBkzEzEFZdp3jFMCTMADQ5EnDyZ3S0s0AO/YkHFTCdFNYfcsGBARIKNL5FZdgIfVKhkMbw0AU64MuCE1bITedGMjiCWA8DznG0SGB4FIOMwDkXn2YUBvgeJhgb7M5o/R6cdO+kTioSk807Id+9LZK4FOucnCibu1RiygG17Ji7j9bUD49sixOdA33x23r3+9vWcAlbt6z8A8dQ9zosHXvh4i7rAwI3v+Ujnwg7CRHAkQZbu+8Yz0osLNlBx7zuoOc/SH9zbgnwH5BGSjx6I9iEEJqckA++2eR9wbgYg74Ea/ovtPmG1690IIERMLMUcucejWdrZw3T6uCCgis5ZMQAvJ+NgNcqceq3cKJ0CJVKQkLwNRis5FmUmZhdndmWhWVZWiOk0KBAjzNIFgtmau2d0xBiEflO2aiMBCkwoLFy1v3jxOh6OU2VjPy/pcL6fqzWp1ej5SkU+hT+2Lb3/608/cyV27du3atWvX91i7Ab1r165du3b9cPUvf/Lf2FRBMYE/2HNjXs5R23ogkDVui1LA2rpeDvOhiJpbhoAz98rMpCTCqiWpFEEsUkTUWvOIAIsIM2+r+WWEiMOdiEQkerLOiMDc8cFmVspELB5EJGb+9PxUa/OAlMLE2TqRQUXL6Xy+rCuLtPDV2vO5ni72vHhzClaZynn1T+f164+ffvX+41fvP3z16fxhqc/pRBKucN1rzzQAr9yqWxFjEDN6rls6iyMVEQFiZrfOcyBOL54j4OZaWFQQYQHz8N6qbvNyKSOHSHSAsJullXz14DaWMYGYYxi5Oaqi4ubWIRXooN3P+HedSlxUx86He5iR89HZT3jQeoHhoPI41bSwZTuBFwa0tebuzNSa1dZkbI8tvu29o1tmgfN1G6iQnC0entzteGGPAgg2M3eXbG9oNmLySNqy1QoGi0REmEVdeZrAskGHEdHT8FlscOsRXTcQ4wU+2B21QgTE8AHf4M/MEoAgCndYg+hmRt+f/KvtPod7/kxut29+G+IfAdu8fI8eGd664WGL+tKVlJLx5Hs8xcujf9e5DnhMbLWZ4ZcHbcZ+HvY6/QKZ6aWOr3GPtZIIi+Deoh2x7twvbaWXu7O5fe2aRE7Hexi8BDPzeDGwAQQ8RIRV8kEQkc1rRneBCR5Is9nMLGsNTjEy768n5DZyrwzoG8++n3s68ek7J1SZeoS5g5URnngN6cFnMMVhPhznQ9rf4YF82q1SRNLQGUGIiXhWPUxTKUWYEV5UDlOZJk0ITGuNiebDXIqqlnku67qcTuda19bM3NbLOassIlqKznNhBhMOh0lEAFdFKXKYp+PxOB8OWqbq/P7D6eNyOTsabI14njC1iEAt9NOf/fy7hmvXrl27du8Bz7AAACAASURBVO3a9T3WbkDv2rVr165dP3T973/wX198rdQqXZZVo4kgjkpvD4fD4cCxsvukaY70/mWt55uJKHJ9uKoKa+J9icXMzdw9OQaS1mESHF4AFgjeARFJoxj8VTM3R4Dc0Zo9n0+1NjPvxhWJ1Rbm4bHWtdZmiNraWtdz9dOlPp8qSIPYI1aLS/NTtVOz5+rvz+v78/Lt5XKq7dKsOnJVOXOyLwBc7V1smcM70cj1dpuLmNNBUxEVISYW0TKnvRoxWjU60qEVSZKJR9AI3oaHD7++Zy0xcsFuBqINCW3ZMcwhIplczeS4D0gCMd9mOIcbd8M22EgDPoK91/dsed8N1TsgComUuDIfiJnchgEd4XalfGxyz2wvJwSZhYe51iPX+S8RA0HjwEEU1n35TrBlJuLunN7fjmzJ2E8rQkohlnBn5jHOlsOb1+zNAXDRK55iXGneV+92f08T3x8usTEeAWHOAXsxsaNTKCghKu5GvaXfS7MyImj0zNsAzC/REy8PP0ocGMnijrPwrVMiiHJKRUCkt8rMloE9xt7N34jw68l/rkaRSxICsFsGBwCgqDJxTqKcNEnQuabBc85lyYHvH3wiIsnJXOsixNIN6JthvvdqRyT8fijuz3lEs+M2PD3YIi+G0YGgwNa3M7Y3D2VOPszdvBdKYpA0XtymV3rhPm9nt11O/p4VOSFiUNrOgeitBZPzDnqY58IiEeTgCEYIkXAWSwLuEc5MRVSYhMFMTGCCgiaWSVUlseNOEQTv60wiPExLOT48mHlr1by22qy1rbomzMIkLGUqWkT65xyr8DTJYZ7AzoxpKhHRHE10aXj/dKrE1WtreP5E8gb2gN163rVr165du37I2g3oXbt27dq1axcA/LM/+Adxepw//odPf/sv1TFzOU764x+9fXx8nGACE7ikAR2ojsFHSBvGOwyBhIgDCYlOOEcQsap0n+TG3UyTFREMiIh5yxwrAAJdlqU18yAzb82XVs06sIHALGprtVqtmUdEeHOvzaq1an5Z7XxeidRB1mw1Xz1qUCOpJE+rfbysHy6Xj0t9Wurz2i4WzQKCCNjIXG48h0GauBms3htsuJXoUA5RERFVZSYp5XB8RMC8JyWJaOABrrYncvl/71oY0sEIL3O+HkFE2fkwEc9uTogkKVszUR1MjxzeoOHyDdszxgp6Ag1/bqBU0N30ZC5HgqRv88gtARed9jDONy9qGNDdTFzrC6MyRhc4N0+KS/ry+c3tbSy9S2E/GdawlvZotnpLVALd5ZEzjC+ZnI/OFIbOcx5usy3Dzd1YOz/E1hWAThMNdxXdNU6kgGSPQRZOE/L2cojAzKNpG7/Gc+eb3APROyvGMCtfvDP6HblCVl7nu29oEdfNYiuQbIZsvyMBRMJVsoeke+SEDMCauXn2gGSWK1OCrpiTFwfcJngg7P7kCFBVIka6++6BEGIR7aeyXfJ9AnqcODFLJtZrXTgd1durvB+NgYDe5vPwd2/2O7LPGGWUzdL/TBUpgdgb+4KIwqOZ5Zbu3j+qmnmz8Ai3u8URv9Z9BkA3Y4jb8715kUGSbKLtwUMvRzAlBpoY9DBNRYQ8yB3uHEERFMEZJQ+AQkUO0yxMQiAhJhKEEm/7ZwDw8BZu1A8RxKyqOk211rWuZpUpoe2ioiwyTWUqRUVUVZV7xY1QlKci8zxli0PAjaSRfDhdTrWtIStZtaX9/f9Hfvn37N2XP/357j7v2rVr165dP2jtBvSuXbt27dq1q+tPfv/314cn0lYkrBiLPj5Mv/WjL754PEY9U1skjIkIbCHRs6h3a+SJxB3mgW1R+Git1m6URrObm5u1lhZYYhbcPX8+WS5Lbc0C1twDw0ghDwd1A7rVaq0VLaIagAEOOGDu1jwC7mSOZW2X2mp60KBz88Xj4nFu8XGp33z89OFUnxZ3RgOsL3+n7cckxyskws13718bq/6ZtJTHN1+AKEOmIGLKDCyyN1wglIVVWLjVBsIIOL8MXUfPMpOq5h9bazFoG2621ircbcXkZrhZgjfSQYZHH/PwbKwXm0d4Y/INAxoRkTzr9AQdYd5zsnf5UAQANw9AVb3ngl+FfLPtYRIwIkQZoG5SE7qnxSSigSv0I1vkBYKZMnsqr4K0AAvJNE1MhAyGp1M/FR44Du/dI4m6FZ6OZCfApEN/mwfP2GeSFpi5tbrWdns5wjxNUwbPW2tpzbXW/Jr7zvRqIIJZMsPeagsE88v4dtz358vzv5tWg1VyP9e2jpXYjObM7RNF9zNzmkWoaDKOzTws+eMiWQaI7kG/sGhfpoVvj3wj7wWosDyWh7CI9DSxd9s9Om39Zu8eTiCREhHhZrXSIHLcj82N9X7jtI/d9AfltoqQIyY3g7a9/y6inpeN4OSRINcZePbWi+hN/BAe7nT1wv8K0/k7howyDZ3tFnk83gQIiIkzQU6AgJWlaGFiYhLmbjQnDCQ8wuFB4RLQgDAVlqIqzMqkIjzWEBCCAFVBwMzCLNwAI3dCiEpRLUXnaQZhqZfE9UxTeXg4PBxnkf60qYqKKAsxMUNEamt1XR+OBxUya63ZWtfz5YT5oQaewZU51vYOp+Oj0+HiX77fic+7du3atWvXrt2A3rVr165du3bd6U9+8l8ttJzi9HZ6O8+TFCkkX755OBYp9cxweLTWw5uenkjarBZmkeQNZkbPQVuEE1PazZFJyS0/y5Thyc30cUR4R0kE4I51reYhRZkFhGqelpG3TrbtuVcWJ1hEbdU8KIJYzHBZ1rV5M3dwC1SPGshfa/Di9FztaalPS326LB9Py8fn1bqX3V2tFyvtu296/b1rC4omyIFFdD5QxhMJzMIiW5/BZubunK3YGGbZHC89OEobdIMkdGeTsOWRe08wdGq2uXcQSIIXIsJ9mOidyrAZxuntxs3QdbdxRFVHXpd6GzQgsmFjgLZ/u2kHIjJzZALaIw3uFxYqU3qenMcUFQJtTA8eMW2P2Bz87cSSDG6WkAGhzeK/DnvCyBmB1logmDpOhJmtmbkNVgooI6DNpCeX+2Xf8xq2+0pAZq+vFYhupQ7wxZb1vnfyx4AH0pAV5mVd3V1YroHYseFnwRe3r72+6tzy+uUYsg1K0Us111Bzv/1ppTL3WsXmP7/I877wu3P/WX64fd23SHAMNIv7xrCOu6TwXc0m98MZDg8Pj6RGv3imYqyz6Du4mtA3J7bNmW24bkAu4/Wx8dg8S2RAdNc7glkiorVMQDuyFWT2dfzOsPNt7ebzf63aPikI3gPLfRJdDegOxKZcRcLCA2Eenr1NKZwQeaIU4EAhnpg7i4OYKaEcJP0QnZWU08C8UYAJLCRMKjyXUoqqainKTOYOhKo8Pj6UUkSotYoI4UGgGW0dAbRmrbW5TCAyt2AO4qWtz+vaRCqkcpRjW87x1Oq//NNffMfQ7dq1a9euXbt+WNoN6F27du3atWvXS/3RT35nkqlIAfGkUh2Hom8nfTMflCnqxZbqrbmbhQWCicLCmq9rc/MAqQhAHnCzQAwO7zDy0jwVTqZEeGSfq8x0mnkzK9NExOGxrq2ZEXM2+lubJRKB0pxkbq2amYo6ooUvtYY7MwkX93g+X1qeZVCLaB4GNMfq4aRG2kgXs+dlff90evfx/M2H89ns0mw1yyX3fhPzzj+iO2E3P0elC9Z90/SLGST5RmZmFlZNoqqwNGtmnhZRdBfOw51FCeTR/U0C3CMZF7iJx17dxL4inj0cAWbqkdQBEEAEBQJETCAmps2MG35lbJcwwpppMjMQtDUWTOBsOFE6hen6UpYWIiIRHAhIYi5uHEDhrrQde9C7QxXy9Ckias6B3qMyLP1BIibKGgWnMfeKpGDeTefWWt6KtIxFxN3N+g0kBIu4e61NE3Vyu5uNF5HJZWJQArLT37ymbhMG3D1uYnc399upsPEfAGLixO8u6zIKM9c3xrinRLSZ4C8d9nTpXzQ5HBDtjaYMIMLSWR07jG000mTOsTWLrQhxE2ZHB3xv/wLXm3hNHd/57NHrKwTqtyZa89bGUN2Oyc3zQoOjcfV5x/tviCLbtvlSjOlyu2sCsiPo3d9p3OGtH5QwLNmbnUZEgMKAAAvCI1xYkZjsGFWnkeC+G/nvzobz/XdvrpkIA9zcRznyCexQ824iXys3mbmGGyIrSd5xHAQiEtDEMo+8M0UwBSM4QihN7c4VyWsJhDCLSik6FZ0mPUyllJyYubCBiamoPjwcA2itrfUS7kLwsAgLDxLOkHiG3ZkVIiiTuV/WZSU34hXeSD58S2+/9Ie3/k9/9uffMVa7du3atWvXrh+cdgN6165du3bt2vV5/bM/+L05ymE9LA8nMDs8TA7kj1NRc1vO3hYnJyYVZXAY6loDzCwJZFjXNT0wETa3pCGn1QpAWEqZRCXcL+ezSilaANTWaq3TPINQ1waQmZ8vJxbVUlYzgESL/v/svc+vLNt13/dda+1d1efe9/g7VCRLdmLDSQAhHoRwDMUeKEAQwIMMPQwQIAEBO/DA/wH/Bs/kiZ0gQgByEsQDA4IHnnnEQGAAJZEZQnCoSJQoke/de8/pqr1+ZLD2rq4+9zzqkSElAdpfPpx7bp/u6upd1ReHn/r2Z7EAMLMUzDKzR5g7iJMZMnOA3ELNd/XrdbMAmJva1uzamgdbUDNq5rv6prFZXI2+//HH3//47fc/ert7NECjM2gf//GY6wck24xuXXgOp3iMIevtYllXKZLDxvKuRaSUOmwDnfUSi7tbBBO5u5ohq9BmiXctkXSSP+5VX2K6rGv2oy0VEjlaL4CInAVZRLIgfbBfHOXac+UW4K6nQG5qcM7EweHu6a+IVHCEjx+z9PLvrYp7atmeMO7ZM0IU7tq0Y3Tp1W9zjUS9d6w/v9Dh0bZmKaUY6DAtLgnoKZADAZ0QJAVJ5cy67/lZOmyXGC7toxWOw8xNeKbJuMe1fSxhQu/bhYTw26mQd88/zcFMpcAsxuBCEMEMo4mO9/fz7iwbYxLDEDbQPgFZUXb086DvTASNbvBd/x1S4Y7opxaIepeZuX/zzBWCocBgAkmejdHR7XGQA0Qo8uxVlFI5PzbhcW67E0vfcRsmFpI8+inCYBEAfhOF8+2c6HFEUPj73PgofOe0zHFmePds9Dr2uVwdtwd/MoY+v7Bx2gGAgAQsfXQmGFGkCDHGWTnodgwKf1TFkdeNsspNfVM5rhBMJKAqsogwgREULsIM99bYfZSsgwFhrrUs6yLCpZRlreta1rUsdSnCxOlpCQ8QpU06tn3b970UIYowU909XKhf/4sIIiZIM+d1NXBDGJEzAnGN+MY3v/M3f+nnvrR++C++/e0Xz9aZmZmZmZmZv5iZAHpmZmZmZmbmE/PPv/pfaW0Ot+b62lgBBwcuwpWLPr0JNIIXJgaRZ1+WiHhdVwBqHggikiJJWShdvAA6ORVmBqLtrUgVKYlWiYiFAzC1nNG3bdes8PUtktBwtgJgJhFRs9bUw1OZrKmgVlfzZrbtquYWMPNddds1gjxYLcxgDjW0oM3psembbf/h0/XNdXtz3d5d96t581CcbNCnz9wPfS7daRHGnc7simtlTv9E/7lIkVJGRXhMIwvKmnefMeieq+ZmIkLMNjrRSYERXROR9z/UCqc9iDRVFBEzNbM0V/T28a34Ofab6Ayg86B2yn5UUCPSf3EYVPJGz8bxWYiQloXbvd7XXPdKb7jFqAmHW861G5u59WfPfya9TBUGl5Jt5Y4ZLe3PHGbJe1MGDRA82ejznXDzfO25jXSbjFK2mxozETOG6gQdsnf2TYl80y8xCq0xljQvIZBwvsAcqZnyBy7FTfNVjKqpweNwRDw/sYiKcOR0yrG1XGmEJ5oFIczDnJiyzZ1l1zzUlFV36n4YInIiRKqKycPVgxBMLLXkKWTRse/9qtFYhTuDMx0Hqvsg7gC0SMkd6MIYdEKO+9x9zoA6Qs+Dm6twbpR7v87RS8F0XrJAKqp7fTdnWuZPIgF03J20dzkVtO++6TvWzRj9m34rgwpLMmjqJe0QEj5EPTcpTqfPEXGc5ATkSZbWjkosfSNgiqxCS5J/BEUshZkQ2oRQhKtw6e4XWmp9uFykSilSiuTJW+QA/ZbqG3eo+t42NfOIWkWIEO5hQOQ/O8mgWRbmReHvtrYDTrSTY9vxWf7+D/R7H22/9Xs/eHEdZ2ZmZmZmZv4iZwLomZmZmZmZmT8hX//qf+HVgeCIBlDALMStcjCFwCR2DjAxk6R/4rJeuNQspRJBqhARM5VSEjoPaUDvkhKBIBFobS+1XtaLuSVUTWST1WYWIRYPUg9306b7vrs7EWqpzXTbtm3b3RzE1+163fZ9a9opC/ZmW1MAZr43Q3AEuyOc3KGOXWO34MuDl9IQf/TmzR999OYHH7/9eGvvml8j0i6dkmjcKospc3jh16q8wx22PlM2GuxcpJRSay1FCKQaDhDlsDsKQMYAwLRQ9N4oUS0FQPLodEEcSocOi+PQLXctcs6BHLybmMndd72bs4eT9iEFIMQc7n4DsqymAI65iG5mOVOyXxLIgYq3qZJp6hjkeqzDjS72ym24EzEiwvUFInk2ORw3iYQp3MvlQtmQNXe3MONSiNjVaDDSRPwvapcBmGZLvpPN1pSJWLiIuPu+q5Q+nK3j43SRMJt7tqdNLVeplMLCfTYgwMzuvu+tlJJj+kwtnSEiIkVSbgD0AnguV++co1vRjzDzsiyBMLOUaZgbgZLjExEJU54SalIEIFPN+nxripx9l8IT5loKEVSN+iUJUtVNlYBSyrKsRPCI1hqG2+HuJH9/cGJvJx9Xm553zYlOWoyAD2/IMcSS05HivaJ7rHOfd3jq1x/7kINNw1M743y3YNFncJp7WPJrujXXn6k23pO8vEymO4hPvQYhJKlxyneIKpc81QBk4zn/mRhXCTqAzg8JUGftB7QnBnFAAEEkyyZYv5iEoDDOUj+IiS6VCxPca+WllnVd11qXWplRS7msaymSUytVm1q7XRUyB4JZWrN9b9u2sUipVQTCXIS5967zX3cplwtIrte2q17NNkRr8aZsr7kUAi70jX/93ZfWamZmZmZmZuYveiaAnpmZmZmZmflU+fo/+NVf+PYf/O3f+K1/9g9+tewtBIT4sMrnPnx1qVKYq4hISVGvuQMsJMTCRIcZOdHb7WPuEWZGRLWWfW/73mK0LN1czVprzBSBXVtypwhW86aaoonEqRGxXlYEVFXVACq17nvbW2tmkRZqFg+YOSjl1DCDG9xz2B5ZQLPp7DDAmHbTzfRp1zfb/tHT9oPHp48et7ePewMaYPEMTb0MoJ+zK3rvu2R+zMeUwpQRMMtlXc8dTwIlrANRekxqrYjQAaBVFWNjqZc1MwTyECDgEdxrpBjd08NXPKQQY9eTISbdzhGC4Z7HK3vrRNx1GRH5ozR/JLRFajTMD2kGmMbovzFfblDAVKYkLi+lUJ+hd3Roj6Vi4rumbULuiGDCcrkApKbRL12wZyWWbpaKOIqud0Xq2/HKZWTuwC73nJiQVfQB7ge1TChOTduNRyfu73XjpKUkTBFQ1QTTAMzMtK9tkeJucRJnew7bJMiYPPn83Or7ABHukpC8qOOey5TdczeLfor1W8wsteRjPRNGRwLoLG6bm7pFQJhLLZ1WDko7fDGn2YyJobvewuk2W5KGFOX5zo+1BbqNhAIUA7QzU35SwN3zNhYW7vqXXhW/PQ08wt3cLSyy3k59mGQ+dX/U0cE/7/h9vfz+7Lrd7f29Z3S9tBdERXRNczJootsJdGwgkDIUz/cfIMyFb1IOjuw+BwEUxABHMCLb0BR2jESsEQtFFVyW8rCsy1IXKULEQiwsRUREhEXG283d3PLzItlszh54rhIH2t7cXGqpdalLJYqlloeHtRQGsJtSKbyuzfG4bU+bNcOu7arRbOW6tbr/xre+99LSzczMzMzMzMwAE0DPzMzMzMzMfPoE8Jt/89/7w1/48Id/9YOnt8LFFy6vLuXDh8vrDz9bhQoiP1e/bzuChAsT5+ffvZscjiF5veCZJdBlqdfrdds2Zkla5O6q1lqrtQD0tG8+fB5mfWBdwsRkf+u6EsgjEAlvxczVEkoFQGVZA5RFSA+Ek7ZQhRs8kCJU91CPvamaWbjBHTCix6Zvt/2j6/7R4/7Dd/u71q5qm7k67PZB+r5E5+XCe+wKd+TtTi8w7NXdMM0sy7pmv9U9y7DspunTCFCAiwh6b9jd3Uy7mGAUfcMNIBniZjNLNOUj3ZkicmuEAkC4BRGJiLnhmBx42A+Gf/o0yy4BX066Q7ank5AOjzH1T/Hfz5E7c/jkw6UUIljaZrPyfCunPq/fdgCNYOJSKxBmFp4vik0tIrpSY5hMDgz5fpk3kfHg+CyJ3WOsEsvJPjJsJBERXfGc097OtdyDbR5nfiJsDAVH3lJKyf76bf0HY5WT9fj8st0j92HsDB/rQUOIkdcFYlxLGLf40IaMZT92d/w9ZRYezsSliI93bJ7Q45qF97Xof883dnjEqDfTwLvvAWgcFfgsAGO4o4+3R95GxxImbR4TO4f1RpjGs4d714S4w46O8wHNx5Zu/pvjNBwibNAnAOixy/1rdp/7QE9GVIoVNMDx8bIwpNi3j0ogGKfXKkR5gYGAXAaOkN6YDkYi6S7iEAIJkxATrcIXoUViKbIui7AUlvzXIB3luZfM5GHaFAiPUNW8xOCmEQ4KSWSdGm/mZV1KERaOcClcl1qKsIgTG9NT25+2fQvfdvfW1NGcm7FHmcbnmZmZmZmZmR+dCaBnZmZmZmZmfrx8/R/9SttJ3a/WXtEDC4ioVH69rg9rhartm+5XAhdZ+0ff1Q5lAQD37m4upbS2R0QpZd+3fW+1LsyUyDUrzq9evWaRd0+PAAnXdb0ApOpSihQppbTW3D1rswhIEQJn7zQC5tFUPeLy6lWAtl33rZk5QNvmbfecUqg5jAvwiLa3tu9tb1vbLIxrVaItYFyuRu92+6M3bz969/S46bXZptHGcMIzicaL1I2OD+5nBu3KrijdHLfpc5BlQbZoLdJA4trCnVikVJaCoSZorSVsfUZUk0SzSG8oa2MWFonDmBvBwmWp50dFhKkRUaohQN0uTURF2CPMxtTBW8m370mRfgkBXfohp5dPCaZpQNjzMx5MXJgDsHCRwizn31fjdBahU/BPPFEpXSUIZtamplpLyf6yqgZQ0qB9/5D8xuxwaveivUhZ1zW14k21lpJoOFXjy7JImpQH8DUzd09fx7HBcykWQDZ8E0Dn/TE48EDeLCJZW3726txdhJl52/eIqKUe1wEO/bS7m1sepojI20e1nGz4LvK5ailpcTkfFCIqRdKenJcibmyZulY5LHoxd2jCETm4MxCG8NRSPzs2x0UJEIEJuR0uSJLuDQiQEN/k0TEuhPjNFC+u5jaMODkH1B03pcxL7LvLLvqI0BgjMY/35yc/5HYPBidEZ/jKfGGmcPTZlff6j/FvgpDwGXDTGKWYrmfKAZEhDulTBKnLPYgry7LUdV3Xy7JUfljKZZFC3mXlTQkQqYHI+aVpKqEwM922fVmWUvIDFvmvYiNyZqqlLqWusrx+eH1ZVy4MuIc1U3X1cC6FSJzx9nq9eqiHuuHj8te//e3v/uIXPvrMq2/81nRuzMzMzMzMzPzJmQB6ZmZmZmZm5ifJr331K3/9Ox//5//y3/xPX/1KWS4G4hAWX1mY6Prmo2h7KbVtGwK1VFN1sxRAH6XOlBGnATk/QV9rTftB9hWJICzMPCTLLFIx9LVpIXD3FBG4u5ppMzXzcIAjoO5N1dwDbAE335uaeRjano1htoDB1T0III5wV1dt27arKQprhHoEi3o8NW+OzeKq/rjpu609Nnu76dtNk0QzYIBjuKHp3p9wZ37oX3qf81b/7A88dBNMhVKqgV6wZObU+CamHKtFcWqyEndFBnrf1lS1lJri5gTH4Y4xWK/7EHCSpBCSqx6gucgJKJ9KvsyUk9z6xs/t3xjWhlsb9GjM4iCuo1p7k2UMVzh1Om1+e9K+LOfRdrftHDt/OC0Sod7k46M0fX4pueQYhpAIMBMG1SVikdKrwKYk0ovM5uE2ZAc0CvGU1d/jqEa39w72mjeNQ8XEvdY7dp26NSWYJSLCtNsdEFk+P+56qD96yTeHEILHi4jehnbLUygi141NWwRAjD418VQTHisKAhPnnvjoIo99DPigzrdjRkQc7iCQSJjDDWH9PjRk5MON3A3JvedOoHF2hXcryzg47h3oR2pGAOrUuxs5evcYAQ+MGYOfZHCmfuvoR59f1yeEQSnZGKMFczAgETyXm7qJ5PnTHX/nPhryeLs7EwsTPLXOKZKOElyJF+ZaCjMx47Jcllqk68cRbsJROPo8SyY3R4ClhKfwPgvg5Kp5makUJkLARfoowlKlVlnqUqUWrsI5dLDlMiqClwXCT61t+95Aat7QNnVs/uGjvv54/+If//HXfvSSzczMzMzMzMyMTAA9MzMzMzMz8xMmgG995ec//uLr/+evfqk02oqBaoSTGwKViLzt+5U8Lssa6uHG3AfuiYiZbdtWa621llICjoj8Pie2pWU4IhKDJoAO4hzglftw8xgQmXtruu17eoc9umnV3JvZtre043qEWbi6tQgnlmKI5rZZCyIukkpcV9tba02doO6JLz3Q1MHFiHfD466Pu77b/QeP+x+/3a4eu1mY7e7J9gLo0oD3Vu/cvX3moyDwnY4ZJFKzSnzYjI9BeYcIN3nzcPWC03cxBMGp4HCzkqt9qCX6mLw4YPeNX/cnutVpw6MrkE8i57y/MOeB6FcXYoguhm36gJvJcHNe4rGBl1Zo+DYCXd9rnlg9nRvoDg0+8DYGxv4U524AkSsTB/8Hhka5A8njRXZw3IuzEabo1wMQ4chBi+//Wv3slkC4EzNyqd3T10wD2qZiBrdxdAPIR1BEleLelgAAIABJREFU3OreNEQZiHR1H7sbkdKVhO75ivLMcWtEgn7RgpnITQMAS3+rdGaegpGx9DeFyHvykwMEiyDd5fBOk8OJiWtNNzNC83LKbUMn70oeiaG/GCZyCiIwUT9v8lMU5jE6v+PtbfeIOc4ujx/NoKO/vNP1ihuYvh268cGEDqAFEHAJJpD0AxljiGEMCH5+wpvxg0GcZmsAACM4jRp9jCEEEMJCZWVZS1nrkm++dVlEuAu2w8KNEExRSpaqaRiu4WZujoiUe4QFE5UqIkwcEbYsZVkqC5XCIiwiTAJn97TKmxSRWk0KiB7362ZqoF2tufvW8Mvfxe9+ET98mMXnmZmZmZmZmR8rE0DPzMzMzMzM/P/N1//bX1F2Z7LiaBQOAl0Irz54YBE2LUAhlvQAsBwa4tZa+gdKKWbqYeuyiJSUJKiqmSUTGlpecce+t6fHa0QQU5Gy7VvbG5I8uVuESFkvl+u2mceyrBFoZk/XDcx1WUupEaTNyJnBTLJZe2rbm+uTEw4CDg8zVbMth+t5LFII5B57s928WbSgBm5RPr7qD95d317b26frm3dv3277k5oNNYd/EgN7PwnB4r3f0Cjbk1kdpQBKLbXWA+UluKQbABvz+uQO+EUEj+pux8HuHqFuZzdxRPA4Tq0198jjBQRzNw9EFlaZTTU32yltQuWTycHNY2g6MAB0Dk7s9eLoDeX3XnWn96nsuEPhB2Qncvfk8GMdXubQzxj3EFN08QUT9bGB4aaGADFJkST3XfbRncthaszcPdfuaVV+ATffP2MEwp2lz1FMDA8Ci5RS2r5HhBTJiwKpv2Ai70MdJS3qLOzmbg5TEEFkbC1EONUfnce7dUtFKYjQ1pgL8opOL873AnJWy0UkD4ibs7CUclZSMFEReWbSSIF7GWKTQFheWiASkaXW3jeHHQsSY6NHGbqfJL1O3YXIGDKP9J+YWdjhaPEw72aPO8NGIPxGzPt2XlBwjDfjQN+3h9yg+9gHKlRyibkLN0Ly+8CYc9gf4PTsOW5KntwZAbpqY7xXGWCCMAlzEanEC8tF6lrLutRaCnmYqpq2tu/bFuHMVNf8V6rUpRCTI1pTba3tu6uFGweEqRSpUtdlWdd1WZdSmTmWpdaluDUzNWvmtu96fdojIFLqw1IfHkopm9mOMOJm2hAe8Xl8/k39nq4f48sff+Mb7y/qzMzMzMzMzMyPygTQMzMzMzMzMz+d/A///X+KzWhrrS6FhYhr4Q8eLp/58DNLBLtlm7HjZ0nW2YW5IjJGmLmf2rOIIKaIaK0BxCRmcDNtQwLLvO97a+3GWEEsUmt993RVs1qqRaiZehAJl8LE7tCm4aAgJm5uV2uP+2Y5sA4Ij/wou5pv2pqamRcWOExN1dWQjzbi5rRpXFtsGlfVp31/t7fHXZ9Ur0031SfV5v7jkOhPKNN2kkwBpLmEBpKmXt/kO9ycjWkmGjKKeD54rt/oETRsxbnyTJyaDx1q6TwgSV0R6C1XFleNCGI5IO0Bf4fvIpD9zFETpl41PVWg39fvEmhMuMuacMpAgDvrNAhufi6C9917H0A/+2u+agRRr/0GIMIRoaoIEHMpki7yw6qc66BmicMxOvg0xBqEm47i+Q4EPFyY0wRtHgf5LbW0fQ93KYWYMNzQ46MA54GH482RTzquJZj3Lbuf+Skwiu2UtDVNLYEuV8k9UUOESOkA2p26J+d2UAiHEGNcSBimb2EZ+2B51LuY43YadjdKDBkLHS3ucTczNwt00h/DppLCE+tHPDUlkYaJQPjYmaN3fKtCn+rPLyTQP58wbqDEwaN/3lXNDCpc8i00LCFBR7067g8z3f48/htd7HQ65zhBZkodB2ota61CJMRFuJBU4sKCcIT17adWmkKYpTAXIenqIYe5W76/CBBmCiegCNdallJrqbUUKYX7LFgbnhgz1/wnLgIMBotcLnW57K6bmzKpRXNvFHJppT2UqA94+Cff/OaL6zkzMzMzMzMz86MzAfTMzMzMzMzMTy3/43/9N4yFC8qiuq8il3WVD169/vzrDwtLtCvcmLkIi3T+ZGoekTQvIq7Xqza1pG9CWeqMHMIWRERmRCBJ+wGACFU1d+6G2WOwFz9dNzVlZjVP+gxmgCPc1JtamIUHiC1C3ZqbRThIW2tNVdUDFrGbNjVtxsRh0F3dKWcEgimIdvMIJhQnMZAirupPTd9s7e11e3Pd3lyvV9MW0TwswiJexNCfqiLdQzfcnL3gzsey30xAyg+CmMDUmeBJgkG3YnQvcR67dEdxjz/u27wRgXAiIpFIAC0l9+uA2zQMId2WEBHcfQbCVIVzmz7QOtNRsCUAQV2qezwpd+sFvdCADroh4ESt96sZHbreGKF7mCkz9eVyN/cy5grmLhWRvP3AzS8B6PBekc5X/VxUca6fm8cBoN3dPAhgkSLSWovwvDiTP+WubO4SirQ829i3Y+OH0iR36Ti4x90SE9dazcwjiHrz+Tar0Cxl0+hc3gkpeBkQdZw292dufk95CNxN1dLq4B5mpqb5uIH4x9eTH+NYLLPeB8/acozzFR63GYHHwbv9X5g4Q+fx0095led2llAQRRowiAGO0XcmCMqt3p4n5iHrju7ZGT+M414MKh3YB/c7BCOEwGBhYiJhuizrw7py93vkfyAg+8xuRqDCwiLLUi8Pi9RCzOptb21r+962MCWPIrIu9dW6CpMw1aUsS11q5bHrZq3p3vbmbjkgsmtlmOuyvH71oTM56GnXDbaFN3Un/cPPf/ezjz9XYuXi3/jX07kxMzMzMzMz85NnAuiZmZmZmZmZn3J+/e//xx/XN9/7wu/8B9/9W6gL1aUyXXh5tS4Mh+4USmEMCPO+N80uZ3iEqZl7tpjTNezZjhUpAIVTBDGxsHi4mbWmQBCRlELoXWlzB9iH6NfNzdLvwESsZuZm5lnjbU3N3SJ/KCB+enra9l3VkmM5sXmiQ4GTa/SBYeAgeERTZZLC1QF17IYQVuInxbu9vdv2x227aruavXvantq+q+0RerMA3Gqcn0zOXvyd7SiS9glvCIhId/66uTsoXRqMIY8O3Ogj88HyQq0vUmFhYTNLznYzPg8Md1h5e2E1ZRHM2QXOex5hIt1bZ4tMYE4AXZiRU/kGue2T6E41aaKc9daBaUSk5/oZgAZu8/wOznma05dbzu2OOvBYitFKx3F7r0OPHH89XlECaLn5QHJE4Y0703MEPTYVcfSacVSnh1P7aDoflerxigjDIn5uYcdJ4U1EcqpCH0/HRCLSD6tIioLTGk0gOyrHABEYhNMkyDijXSA8LwLdn6HhWY1ODB9uREwsYAp31wYSogjXMXpxrIx7d10cS5VijdErPpb+7psTBj4fn/t8IoC+neunynR2pfO/QrJK4eHWYATFrck9iuXRC95jC4SjOn3blBCvUpmIwo/GdC2lCDNBhIVZmApLIQ6zMPNmkX37sMKllLIsS62lFFmWBYTWtn3f97artmBAOK+RXGpZl3qpy6UugAX8UDxvT1dXJZBqa9paa7XWdVm5sJQiy8JFiApD3un2pKaEq5mHf4TrUszr/vjw8b/6V++v5czMzMzMzMzMj5cJoGdmZmZmZmZ++vna1/DFj//Sq/0zH+6vrrwSFQaEZWU8rOvCjus7Dq8sTd0DLOLezNTcLMi893pT30BEUmo4+rhBZmZp2tJgAICFa605g6upprO5GzpY0uHcPQ4saZXdWysiIkKjLJxEk1hUtTVN9UQAwaLmZs4kCIazd2dxeIR1nTEJsQfUoxnAqebApr6ZNbXdfHd/3PanvT3u7bG1a2vNfDdr5hpQpCj3OTxLsnn7rP9oLXc6GYOqjd/peHgVklASmJiZGMJ9TfvXxMPA4II5FTBRJhFnfbUXrLMpetC/nN12INFBdzs5PWwhue3oAxBH1xS5RR4vKF9GdAXwuFN/rYeqmChuxe3bxnj0jW/OFgzGTjTqsdRtEreVTaH27cWPLTyDm8dww0MAjWHSYOIk3Dn18awPPl4oaIxHHDQ3QAfQ77vclSae5e7hf45BmW8d4QGfx1y+4wW75wWYTqVV07uS/VkmPo5TzjnEKD4PoHzMBaRRcKa4VeLHH5FF6fv3OWGQ5RwJ6OOYdfcKSIgAt2yz9xM3EK59TWg8y/BI4H4ZP0We8f4zgH6Oqk/FaUg/e24MWogXEQ7AgwKAHwfu7hDE8a4DgbrZOYcKdrcGCctalxw5mOvBRPnhhETVwNi+g8I5shnNwszCTCLcG+oEMHOE7W1TVQ8nglQpSyllWZduhBYmCrirefOw1Nu37UoeVcphb1nXy3p5gDCvK0ppqo/Xqzq1sD2s7c1b4Le/2/7yFx4/V3/jW9/7cQ7EzMzMzMzMzMwnZgLomZmZmZmZmZ9Vvv7VryjJzuvH5YMPtx8ykQSthV5Vfl2EdVsI5gxwXapqa7qrazM0o0h2Ew4EMViqmatakBALsVyv14i4XC4AmKnWJSJUNSLUdNsbEZhlWRdTV7OE0cwS7ntr1+vTsqyXy+VyuRCRu7WmHiCRdNqquqezANSatqYIAoSomLmZq6uqq5q6JRLNGqg6ImABc/cgBwXIQRZojk3t3b59/O7x7dP13ba/29q7vV0DW8Q26p4eN1BKQE6iu7FZulHI0+Cz7G0etLJTtRRwACmDZmamIiwMohgYbAAyvvWWATUF6KjrJkFOYHr0cFMT3TloQuYIpm5ywJgWKCJMZKMfTZSY1fqjxj1d7WZp6LvGJ3A8eHVELzffmqlxr2JAkvVwT6ZJOU+vm6gDQBqrI4KFZRTGzZy6eqFv9rzqGNQYdJDIcctAts/xbBdne6SyGcQHCh9xAPBwYykAuRvRqb192lTCy/Bw8whPfwIBYQqApPRT0JRL4VJMW798IwJwuMMNCNSaIBjhFGNGX7ofuiDjWARQxG2O3/tYWAR8kp10xg7KU0f6ucKgGOeHm7t7uHWDc/SrGQm8+dPqM45LBXGc4XfLdfPH3N4gdL/hhUthGXcOjHmA5P28ROQ6d3I9PmXQvz+8GQISpL4DhaiIMFhE6iL58knAzMISZnBHuFnON1Vzc49KtNT6cHl4WC8P6+WyXtxDtW3XJ227qmpr7gqKmgXmy7IstVZZ1stSahXxCDPbtk2tqe7NNlAIE7uvIg/LWiRHvZZlfajrxVmupm+eru9su2rsZuYb3i2//J3v/M6XPvMugD/6eA4anJmZmZmZmfkpZgLomZmZmZmZmZ9t/vE//LuLXmvYhZxag7CbXzgupay1tq2FNWEmWIS21tTJUGqtwiwIomDmUmp6MMqyEkviPmautWQRdlmWAMKdiMx833cWEeFSCrK/6ZFYjIjMbNv3/Hh94lEA1+2qau596BcC+763pkS8N9225hZmoeYB9ghV29MWbWNyIiHyU/vg6HKGyFlz5mGBIFZg99jNdvPNkf89Nn3c9bG1ZrapXZv6icJG4uZbh7P3NoG4zVobBdPbVxAipROdnlHH0ePr2Bp6aZWHNIOJiKUD+4Ronurq6PqGXuNNFO4J6xygdD4gGXqcxRFDAzxwNRLvpcrDU9jQXkC4o8n6PmTsvVyKXis9PTZROA1Dh5lGpAGkb7DT5UhlxLkwTsPE63nb0I50EBkJZ8/ybESqRI4Je2PfceoUp3TiLOo4H7aAB3WHhh/bP60CM0uEhfuxqv1mFnfL8yDPgL5nlLscCGIpx8bzeOQhScE6EU6YvY98zFbw0LuAX9rzPMoDTh9XAPpqEHJeZTahPSzni1quM+DD7BxHxzoBND4tgz6WuRPv8y0Hv0/N8/Bj3JWghVjA6ADaCcFEOcax1787E082T0O1ngptSmkJgzjAQCEkCxbpL5s5T/3wrvwxChAiPLKeLCwiXESWWotIEQ5Hf0tY/zQIECyUwoxaZVnXulSWPGbpaYGb7ftuZsQEeCBYUKostSzMlUWYS6ksJUCyPgTJ0359NNvc9mZ7aztv8sf0yvfXT+3LP/jB1z714s/MzMzMzMzMfMpMAD0zMzMzMzPzp5Ff//t/5y//mz/4O//yt3/9v/tbTk4eQEhwEV6X9dVlrRzsu6l6sFMppRbhQiAEEUSKmqtZXS7EZO7ZCRWR5HGllCxZCrO7t9bSwFFqISIEUqmBAIjcvanmDMLkbu6+J29Wi0H59n1XtQ6g90Ykan7d9iyGmntTUzXzzlKjD+dDgA7vQkS4ufU7kAEGGMgABSukgTf1a7Nrs81sU33cWqo5djMLtwjrxO4AlsBwDdxC732ftc7oAPo2Ig0nb8FpnB3xUYLmIsKS/DmxVn+BoOTTdDgpIig8vEM3Zuaunrih0jRJdEmxRx+jly8lK9ARHupxe2WZGAB6YFUaPpC+2gEMAH2Km3V/iAgB2tpQRqfwAmlPpmGgGM826tEsoK4OSV7r2R0GUnB892Qx1CH3ALpfKYg4nCmnh/Sf3neHT498JpUg6qDZnXDMGCSAkA10HM3x3kl3d+IsfUNKSfeDo5/aw20ymOoomB8XAKJf3OhXKThe1lpb9OsuYyUQ4b1bPfY9IsIt3MOiL+PAzbeXPZ72/nLKJ+X5WX8C0DRY87g9LTO9yg3gzp4xquaeeDrtGRQxxgkGA4LeihfmvDqRp//pmg0YVAhFijAT5ennEZ74nszhHvByvKOEi0hJX3uqcRCIsBxMmQQ8IMylSF1qlVKKCDMXIaYId1XT5uFubm6qDYSl1lKkP6SIFCncWXx9+IBk2dUet+vm2Dma2t4cvL+TfXlitOAn+sZ356TBmZmZmZmZmZ9JJoCemZmZmZmZ+VNKAN/6T/4SgL/xv/3u//zVr2zBblSYX6/Llz/3+vOf/ezlcqkUADtKRDBRZQqz9BJs27btuxT2CG06LARkqq4WgKmqKkvpQHnbCXh49RAR2UHsn3zPfqEaqBAXYt62fdv3iNDW9n0vpUZg33bvvJp31V3t1avXHnj37sk7WqUxrow8YBHh41ly/h9JdoUBgMgRzZqZWUADBpiTgx0MroA4uAG7+1X13dbeXrc3T0/X1nb3HVAgpdQ+hrcRTgaOzPu/2R0wLWGYx8u//SUiznJ03psEg7KNo0d9I8f0wqMgi5uS4sS+h4gjIgDmkj9wNxCYOQ0ewtIdICzv7dpNgpFhZiFOtO2HFaT3XE/n2bB/JGPt/fdAwvHciQiwcJxq2kSkqgBEJFG5miViNLNsf6dW4tnK3XrAftsNouPI3z0k2+B0KFC6Phr9Ysgd3b4h2rzYkMRURIQlgtzsuBJDxLmTRYq55bRDAG4hpeRBDMBHl/28vnQj2Lfbe0V9SEvyL/cV73E+nOLmZsbwfnmgX5M5/ffSq/uTc3uW8ai4/YSAPAnH9725LGBhyYp7tvSP8+Q4X9LjnW8SAcrg1wxiOgB0/pX6V2ZmISISYeE+z5MIEWauTVV3taYRDBRgZbmUerksl2Vdl6X06wGIcDe1ptfrY2u7Wyu11Fovy1JKrbWsl3Vd1loXijCz1vY9P3Fhpq3ZvocbEaRwWUpdylLLq8vl1fqwLBcCzE316mFB7OXhan61aIg9vLVmTT//8MWP/aMdW2P759/8fz/tsZiZmZmZmZmZ+fEzAfTMzMzMzMzMn2oC+N+/8vO/+/Mf/ttf+PAV4Ea1rstSHx7Wz37wQS1rqJqpAIIoiHBNE8K+t33fDwKYrLDWmhMDAST3rbWmF2LbrmYmXcERABI8Z1HVPJqGO9ENgLKZ5XBCYkbAItzRRQ/EUqoH9mbuls1PD+T0whQce6A7JQJu0ZpFADHKtOEW5m7u0HBzmNPebG/OUkASIbt789gRm8WmdjW7mm1qW8Rutqk2NTU/3LQ+lvSu3Xy33NS/nrjwXQl66Hd7kRQ8NpLiARqwLLpwg7rHpPPohNbEo5/8wu+WvSF81FupF8RHibQ3qtPFfMdqxz6f1NY0vh7sko5neP9Uy1sTxR7WEgylBzOnAATowwHNDEAtFRQepk2f7VLfLb7ddKa257041piOWXIYqDxnDCb4TDjPbGYIsJztzx22ppIhYTrxWI7IqY8hwiByDzdL5u6Rwzqzpw/pFL6fhDj01tF76nRA3VuZur+yGzHu6oxn8XjOlPNMCnj4cWodPfjjMJzu/2MmTmfSWTnTT4x0ZVTioX/Ogneace4eyMR8czoHR0i/ZJQwm3KiYCEWAufQwn4upEhjfO4hYXb3fUd4MIKFS61VZBG+lLqWspTSl9HcTFXVTcMdHiJUCpcitRYpzMSSKczEIOjeWmut7fmZjSJFQAJellJqKVWCgghZwGZipgJiMMnDEhTX6/7OdDPsaldH+HXbLq8qKvNDffVPvvnNH/8ozMzMzMzMzMz8eCl/1jswMzMzMzMz8xcrBOCbv/drX/2FCrytb773C7/97//+r0Db/tbePu0MWurKRBVOtnHbEYYIgNXM1PID7MKSko1lXVXVTNMtm8SrTxF0V7OmhkSkIil9ZmIQMSjIzYJApdZaq4iER5I+FhYRDyTjYyksxTwswg6NLZGZq7l7qJm6pqHXIxBk5tvWEhV7x9NubhYe5mquHh4sIPZGQkNfYBTpvOZLkQ9Au8emtnlsqte2b7tuqs1d3VvXKHcV7yHoGKuc3wxP9DPuR7iRwePWAOAD03ly2u5YSDVwNzaEJ1LNVijSrp1TI+m5r7mXQ8k7LU+GOrikI8gB8t7OHj6Q8diTW4EwmCjfSPfZb/GMZqa62ofDg2i4oQGAiYmHIcXHbiZQ77qPgzby8EQnVgVuL5HSFe2HFuNewXFah8TB3v0scPeg/vwp6ui1bnv2KgaAVoMEEZN3UTCOAX4AEJqt+4i+vMm4A+ah3ZQSadvu+Pp4PG7o/EaTYyDoo2Icz08XAHA7I+q8VtDlKt5lNC/lJ+DOuZodIvM4BM/k3/l5BAFJ948kQff8qAD3dnM/qQqRkBBGhz9CCMzJnTFOBggxEwb2JxClJN7d3MzdjxdJTMJSiiylLLUsy1JFSuHKIkTMZE1NmzVVbabmYRQhRGtd13VdL0vq6N0jx4XC3ULNbN83NY1wYi5SapGlLGvJGYTCQrvu7lakuHsLMIikgvC0abO9Ea7u16ZPoY/+9OCvRPSxlf/1//o/frIDMTMzMzMzMzPz42Y2oGdmZmZmZmb+zPK1r+Fzb3/xg3df/sz3/9q7f+cPhRTBbqiCD5ZFdLd3PyQ4At4/B3+GhCBmKSXB3QG1SilZIGyt2VAoEFMpNbGOiDAJiJkEyNIrgRIjgtIoTGN0XqQbgYLIzJtaU83Kallqa9aaNrVddVd1s+H6cDNX9bQ7RAfTfnyCvu1NLaQsHqSeZJDCsZs38wYYKF+yeTRzB2vEbva0t+uuV7Mn3Z5sa+7NfFdvAXuGP8+V508mfgfYPd92/ysinW6+gVdENjVrh8E0dN0dDvb79YGFA3oTkQ8efpDlzjbpXpSc9xmT7bpbwdzdaylEZEMl8X7tupsjfPBT5rQen1Alcl6iu5s5AGEW4ehN3xBmAGbGIkUkq67dR0Fg4nQJM5GaaTMpwnSWOvdTtVfliYTJPVprQkwgc8vliu7Q4O68uKsd3/48lhWAo2uXOyYl4BBeHIsRncu/d5Hh1B4/P8/9yqcnxIfJGyd18nljvfN7247f7vTCJYHbk51Pz0OG8d5xjNOMQxykWECciJk4hcgBP15Nms4DLslhwTyejhGCXtePiEVqlULIynCenDEYd5b0uys8e9yWfD+fBYFIQQcVFiYWomUpl3V59fCwLIsIW2v5zm7bVU3dnSwY/cSrpdRahEmI0smR/0SEA5E15ry0k4vgpfJ6WUpdRNjMi5TK1SPL1Pvj9ckj6uXCpXKpRuIOQyhh91BvLfSj9u4/+9b3vv1XvvAHn62/8a3vvXRoZmZmZmZmZmZ+VpkAemZmZmZmZubPOF//e39vf/WO1mt9/fT4jpglwiSohl5qWZZK2tyilFJLIQITj/lpAMgHt6u11lrTokDMGDhPirCID9KXjg5TB+CO5I8AvDdhqfuFEzimUAMEkLmr2t60I8taVV3VLKKp7bp7585ZjAxTD1B++j/3JE0dqmYWZhFEHuSBBM2qqg51aMBBDuIbgCYLMo/NLP+7erta29w21a1ZM28eDvRCdLj3DvNzDPgp2qcv0WcMycH5ZyRpdh6l2vzuhEFBffQf8bGR6HD2pk+I2/bvE3j2k+hm58608zDF85fUIe4dC+3mjfOrGfP6wpGVaKL+BIOVB/pcRgwyfPg7EgELS4rFcyrj2R7S18RjaEAoIkxNRNLXjM6R75Z1oODnL4kikCIR82DK798n78/91O+13J/nLMd4XoePoweNw19B94+ME+Ie+o6XnuD5jS8B6Bf8LdTvfIgySIAkyzzEJgeAPvW1iTp9RnbXBVSEBcQIHpdcCnGqsSnGE3UXyW2YaADhfhwTIip5NjMX5oWlshTiIlJLIQphKqNcb9bMTM1UN49g4bUsSynMXCSvhRHCwy1HF443EBOXvP7FAmZiIRFiJhYEwt1VlcAMthx3CARBlrU+vLKgfdcdBiqWuuftaoL/5Td/57/8dz/zS2G/9L13X/tRJ8TMzMzMzMzMzM8kE0DPzMzMzMzM/LnI1//Rr7QdO+obfv3Fx4+MFKAaWKt88PC61vXhsl6qMFyYRCQLs0O+HB5+WS+Xy2XbtmTQTISAu0mtXGS7bu7ORHVZImLfNtWsKnek6IO4HZMEe585ImuSFqFmrVlru5kTFzU3d2I296bNLCcmmgHuYZp0jrpdw8EiQKgagt2xm7rDQUxi7tu+eYgHaZ80SNQBtLnDAw5qERrRInb4HraZbqq72q7WzNWhHurR3DRCI86mjbME931q+1Jeqr0+u8OJI48nuU8QSyGRu4cR0WimEsafz/wbLwHWsfPGREXEcgzfIdYYSfLOkvZqmHv22Pl+784Ch6wUuzdEgDnVHYnXDz9Xgj3oAAAgAElEQVTFDRkTRTgBzCXcw/X5Qr2/HtyNG1wqMZtpPjOxdNoJIKHj+9A4AuEkBUC0HSKQwkS3tnR6Tl5cq+et4v4/Glu+taHPTxoR8NvYwM7E7+7RB/l9gn/79Ppf+PGLAPrZfZiojJGYXdYcKAEB0SHEABAWsPM5I2AhGWZmIoKAl1LSy9GHcsbputDoOPfuMwCEw28tfXSHTxFZShEpVcpS6iqlClNEAmhTNd2t7dY0J226mZsFeSllWS+vXz0sdaG+vm5mps1NuTvokeJnqUu+L6RQKSxFSuEIa+2673vTpqp9f5moVFouy3qhWpv6FtECao6wR9q/8AP5Z7/zO//Rz30OhP/z93/4I47TzMzMzMzMzMzPNBNAz8zMzMzMzPw5yj/+h3/3oV3FjBrjchV1plqEPrxcvvS5L3zw6iHaFtbCNclVzpfzCDfLsWepgyCC7s3NiRkEj+heDI9AmHnbW7JLd2BIfsMj74BBJCNCXbM67SAzV9UBxHhvbW8aw2LhDvdwtwB5wCySaAXCHeGQUtzj+nSNAMBBef8uagjE3qJZmHPiZhCbe7OUR0cABrIIi7BwhVuERqiHOTRgQPNIKcfu3ix2y751L0T7ea1f/DXwR3Pp9yuqz4vFz0vSAIYqOm+4CT0o0rXLXXlwVn2AAHAR5mcbJ2JyM1CIyCC3z3fLI2icG9lnT0R7A9Bxxp55+LxrkYGcRujuRHynGL51dynnUErpvJjuC9DPXv/5KYsIEWn29CnbugcH/qQpjhEeUgoQbdu5iIiMl9Z3mDn32e4f+dytMWD6rfV84HU63zMBNHAC0HiBQY/DT5983rxMoN/Ls+UjgIlqzqUcP6UAh3PgGNTINy8HhFhS5M3Meajzn4MUQ4sk9XXvpeHDxYHbaRT5vDl+kAAmMHEREZal1lpKLbXWUkTQ373WWnPVML3fFEqRJMvLUtZ1XS8riMzser02a+7KYGHKy2mFWYSJgpikFBFmZiCl9Arvqg1HEIFFhFlElsvD+sGHGni77btTC9bQXbVRbG/Lq2q/9/Gbx3f6mz+c6HlmZmZmZmbmzzgTQM/MzMzMzMz8ucs//W9+FUUD2ri9soVKWYReLZfXl4fLwwPg9vjWdYNrR7/hBDTV1pqI5NQ43VtWnmOYiyPcLFSbezCL2+g+MjMziHJQYCKsY/RcB9DCAfIIM6ecUchlb21v7Zgb1yuVjiDcAeiICHiAScx835ube4CYIsg9bCiLm7oqzNmCHAQmc2/5Yf7wlNJaRI4+84AjLKAeFmQBDTT33bxZNPPm/mRZjtZmpukUSZ9x3NqefefxKUjhy785/km/TxK/d5/hPCAi8LOW7tFtzeFt5x9kU9TdAsFEIE5IiMGs3+fh/aHUp+ON4m3S5mN4IDzc3Q8IelIxd+tG3jGol6ZVLSJKkZR0vLQOw6hAAND90b3yHWbOzCxyLwtBx6bPNhTh3rXUqprnJk72EQKIIj8McLcDcX9cz/w97u4x7MZxuuPR+37+4OObl64/vJBPA6CZSIhxWgsGyeHZAQjBAY5g5PEmBjFRIRai4eXoB+J42x1P3o+bu3d1eOSRS9vzcToyUISLSBEpxN3RzCIihUXSv0EEwMzc1HI0qlm4p1ejCIuwMNeSj+JSRESYuVnbVbe2hxsoikjNJyrCzMLw8AgnCqJ+7SPC3YyJgDA3cB90uKxrvbwikq21R7fdaVO/elh4eYNf/s53/u9f/PL3L5/5F9/+9qdY+5mZmZmZmZmZn3kmgJ6ZmZmZmZn5c5pf++pXqst+efv7X/qt//Df/u0QBtjh7FaJKAy6e7u6KYUtpajZ3vakx0LU/bQRXIrU0qfERVyvT8zy4YcfupE5IUW/IsQcATNnImEWFmYOCjMDg0VyqptZELNIXdfVzFvTZjpMv12WG5Sl7GziUlJpD7h19LvvTc2YOMAevXLbWnMnczYnC8pSsIU3s91Ms7rp7u5mlizTPNRD3dWjeTSLNv6qHi1ic2xm19a2bdu1Jc5WMwMswk711k/ZVL2ls773f5l8wcLxAoB+7oZ48Smek2liZpHE9TCjUkkEwcdFhtQoSBHq4yWRFw9eGFQYYWrcq6ZwdzdnISDcPIcK9iGSvRXLzFlYDvMwNQ+vtbII8cmGcdo+ABHJs856hR1d7eJeSy21qEbaQvoumZ+xad+Uxz1ZBiKgOpQdQDisgfluxVLr8V4Jevz0+OO5wOSlvH92xIvH9dPn2QOFpbAcVwjyWFLk26ADaEIIKIcQMgszC3EVqczkfYZfvkXMfUic+7qdRxH2ZwRz7+GTEBPATMxUiyy1rstSS6ksjD45EJ7WDNOm2pq27TgoIlJKLaUstVwuS8kwFREmDtfW2rbvm+4aTsxLLUvt3JmJas2mvzVVa2q6uxvgIAiRsDw8XEpZgiiEwExcQLxre1Tdg3dgd20UX8KXPt7fvPrjH14e25d/8IOv/aSHZmZmZmZmZmbmp54JoGdmZmZmZmb+XOdrX8MXP/qlZf8Q7eHBJXYyhIcvJGvFKqUgJFrO9hIpwyqcQDAND9TrkYQINN0Ly+tXr8PJLFpTiwDxsq5E5GFuBoewFCnMbNG1BpHzzsxLXZg5QbCamXukUiJH2FlY8kzrAPMA0Kamzdqu3ZrAJZG3e+j/x97b/NiWXud9z1rrffepuvc2KcsU9eUYiqJJBNhIIAQaxAMCAZJJBploZBgQMhAQA/kf+m/wIIAIBBKE2ANxlgDJ0Jxl1LAjBYSTKDahSKQ+SEndza46e79rrSeD9e5z6350s2lRlLr1/njZt26dffbH2acKhed96rfcj/0g1JNjZCQoomoURObh4RlBRrIs0wkEMCKPyqyCkSQ0ACcjEWQkDuZRFunZ8LRgjvDdY9a3k545Ml8VdJzFU74eT978GC/rr685Hp7Wefn0ebdPv7Uv/Ck47SqcLWSeco9bgRWnkGLm/vN51V4WgC/71HJrNd8UGaTUoD9yDrjLSuhnDVtmtRYsY0fJRURYqx14SwB9m7Z4S6hv0wxVRUTfjK3fOoTwlc1Ys/ee3K5SjN+q4+dzbtu/5bXk7a/Xo/O33Zjk29ca3nqDXx5Wnjwqp2FE5HQ63zaQ827gbGeTCghhorUaJAIltKYLTvScD5lzYGgZdMApgAbrlks5OqBttvFJsFvvZmpiVqtNlSO3eYfr/ZSIMZDTrcEkM81UBQJaBc31dFMTNdNmJqf6pezeWXYOkZLRq5opTCGKDHcfIkjG8ENEVbSpdtNuCubL8Z5qoq09exEiD9f9muGgE3Hk7uPB9D/73d//o5//2fw7P/XV9957yw1cLBaLxWKx+GtlBdCLxWKxWCw+A/z6r/1SoyTi8e7Ddz58wehiENE74gvP71+8eG6gmbbWRQRIyZiCXbkVY6chI2Ko6v12B0pEHsMrurXeRAXI8EBSMX/jvpwVIDMZmRl5d3cnqvt1Hz4iQqatlZmRkTUXMZjhp5wjy5eADPrh1+uhUr+V30rBkZHDYxwHRTMxhvt0dJioEBieXhkxkUlnOrMqz16S6NKJQBJISpBJBEvEQSehImZqvSrVu8d+jGMcVZc+mLd0u3J2kakFzqm2xanGnj89nlFs/YOv/FD5ivT4DX6Q4uxpzHjrA+e5nGXqCogBQN44RFmEXwmgRc3w2nZPhvlxdocFlJsfmXi9uv3SYfH6KX6KTnllzXztc9/nWefwv1t5+fzvp+fl7eIZ1J9h/cdEyQDfkkDzY59VCbDUqoecBmfUTRM7M+jbNZ1Bq9xkINN9MbvnJoAklecSiMw/kRHhOXXuSVABg4qIASqoxvSm1kQ71MqsQza1ZqqGWW6X6bc4l3gCAiTG4ciaPTnfuHdb772pSi8htOpc4DhfRuKmukmAUkMxRS739713gQIBBNM9PGKoSjJHjNZ6b32z3lWbipRnRiVV0bYRPCKPjJ04Ijw5PB7HY2uXL3xw7bv/7J+8/+4P8CZYLBaLxWKx+NGxAujFYrFYLBafGf7Zf/8L276Ndv3ul//tf/D7/6mFqel92965u7x4/kz7Jqrd1EDJYdZExMNLkuARycx0jwGiW0MCZAShRtHrsSdZvVShCJGREcGcrdVkRmRG3N/fq9q+79f96u739/eRsR/Xm12h8mqPwCy9VgmaIsbkcTiTpAhU1UwtKZ7p7qYGaETuxzjGwDlULQnWhDIoIQEeEXtEohJ2TUgm3COImxs6E8PDo8JrJpCipeyYFWlmJFMEqiPicN+PMcYYHgCSkjN4L28un46lq8b021PP1+wcb0miP5WCQ54E0J90oDcf04/b+WuZp8hr+fNrswQ5T/XUS+PNcXtzzORbcuNPEwrzU20obwuFiar6nrvINzb5NLxy7E9YGXjrOT5tMb+e95e2AlSR3ppWml+18QqR5dXLIoScsyIhCrZmd9sFRKmRGYFaYyEUAp0K8ciIU21DkEiFNGmm2k5DdFe72y6btibWW7l1wPRMJ6JMy8kI93CHzBUXM1NTQFWszM5Vdr6/bN0amKIzW2edw1yA8mQKpHVrTVrTbbsk83q99m1TVSYzjogjfIiitbbdXVpvUNlab9oMGodHuIm03qR1afYwjg/2Y0BD1GNE+J893P9vv/d7v/yzP/aTL9r//H9959/r7i8Wi8VisVj8iFgB9GKxWCwWi88Y776LL7z/U5frF1q8013utVnrJmrd7u+ePXv+rDF7HumeMzGOzBQV1Zr7lxnhYyAoFNWWgCdHeAJVMBWK3KayCSKmdllF1MxUK/k6jsM9emsEPaOcsCXXeKr9BYSJzBSxStjS0yN9hFnvvScRmR5u2kj4qAI01AxQAmN41NRCKEUSHORgpczMCp2JJOZnwIqPIzKCkfQMTwZ5C6ArVvaISCbTIz3i8BmiV1qYiapxBulg1AjESuzmx8kzneSbcebto4/pML/K6xs9zUP55kZ/2R9j3xK3ypvVaWAG0G89xVmI5iuz/j5221cPftusXrVTU803s+yXbo2n5zb9yJ8uw/6E0/o+/o03k+XbZ+xsjL+MoadI4zYWMqWS6CnWyNtpn1aU2ilr5GAF0Aat1RZTRZ7icybJ+noQnC6P2d9OFdHSQquYShPTajaLluK5W1MoOGNxIcfYw3dInlfE0kyLQFTUtLVm1rSGReocLWiqzayU0KfxvQaPnhE7E6AK1MxMVAVT4p1zRmm4gKbSmvatb1tXMxIeUafatKmYmKm2q4/rcYTBoXvGEZ4i8uC/9W/+8D/+0hdH2u/92Z99yvu+WCwWi8Vi8dfICqAXi8VisVh8Jvn1X/slTTQ2xP0drnlRiJlaa/rO/f07l8u4PhyPD+G+71f3o6Z+mamqpvv18RGRQmmt1wQ/MSHhVesV1RkWS1mYM0JVW2vbtuVp6q2hZABQPl9QRcyaqgCICN7SwQSThJjZtl3c4zhiDDdtrfUkPcLDVYzEGEfF2K01QDK578M9UHJZIAkHHPCkR3pNxCMISU5nCImkRGQmkuLhHnFEzOg5GWQmPSLqsYxIRuV8JCE1xy0qgAYq8h7JzCkaCWZklBiEczPmmzH0G86Nj8lKX+/wvlXs8MMLoD9O7fFGKv1qDv5xYpFPs/dXdvrqhrcxiW8JoD/m3J78+wcLoD/lpvLqf/Uslt+O28Q+IYCeR5v9/5dHroflfFLFvlVVLhV0zQYESmKRKLU6CEEX1XmA6eDQOalPmrVu1mp4qGgNMLxpP1SUicgokzOQ7nvEoUJTUTUFm2nvVotMrVtvzVqrlnP1tW+qjTKKzMAZKZWqa10PVSBajm8BOMYAUk0zo/400633y+VyuWy9dwI+/LofEGmt393dA5qej2N/zBzMAWTEzjiey3aV/++7D+8/HP/Hdz78lHd8sVgsFovF4q+dFUAvFovFYrH4DPMbv/qVBr/c4yd+sn37Dx5VJaSJtM2IkSIYY/f9gO9bF0Eic9uaQjJCSEYOD1G1tl3u7oO8Xvd+ufR+aa3XhMARrmbbtm29V6fRVAEMHyKqqiBfzkUDcs6o43RAT0nvDIUh2lobwyPYrJMSkZE5hu/HISJl+3CPyBRTERVoRESUVhZ51plH5kh6RkR40COGZ/WgeU5kGx5MUTXP8MjDg0RCSnhAMGOGe1mCkswkk6JqBCLn6MUAhmAQIxkZGTEykgnAIyMyMwMMcDCDeBpDvy1Efkskzb8BAbTIGzvl6/3tH1C3/Gm5da8/zuf8CX6Mvzpeps8ya8Xy5CHTGUDPhRGgliduT51BM6G3MYMigNg5cXCGuTPDJcp386RPf/ad59DBy7Y1q4BXFBCRbq2bVXNZIWc6TEYys764kqkwYs54JBPIfmm9q5ViQ1UEremlNxVRkxpIWLNGp1nDvXZnWnMC57WTMadWTh93AhRFM6svxPJ0CNi33lubrWzIHCOpompJeKRaF7OMPJhOCWaQh2c6t/vjSjkEscnX/vc/+JG+CRaLxWKxWCz+0qwAerFYLBaLxWeef/nuVz78YAjw4gv997/1oXIz6JGRHgzcNb2/tEsziZ3plTFlxDRpRKqqWbO+VRDcts1alylcxuEDgKreXS4qmpmqBqkYC3Ns2hkPPtUFEJjZMBEZ4YkyOosOj4y01t2jwujqHbt7ZqpqVSU9onrNEZmVFyci6aw5h0xIbQaIJ4/hok1Up4c6OUYkITAASY4qRGNOert5QgTgbEafETbqsuSUe9ClRqchSWYGk4CqDM+oFFslVY6II2JE1N5mAFjBH0gigYAEIGduKQBEeIsH5119qyVaPiaAfou04lU+2Txxe9rrumV52/M+oQT95Pk/YEz95HlvfeYn/tT+0mXxaY7wGnqG3y8F2BUbz7mDUjlyUxWIVqmfJHkb2VjJOYD53joNG7OnXPuXUprf7BxzGUQ402c909u69SpiqgpRzjGBatq2riKcb18ooKoqUikwklPxUZ5oMvPUpJ+l7NZauZ0vl771JqQKRIRIVWlWp1axtwIYY36BzKWZSAFV0EybiarU9E8AzVpTVZM5z9A0mWTOr3mT+n9Jo0sKr2Zt26RtSdn3sY/jAEXFSU8Cfjz447/5w2c//+X24mI9vvretz7pXbBYLBaLxWLxN5UVQC8Wi8Visfic8C/f/cr7H+5j4PqR89i13Q8iIZvg+aYv7i7P7u9b06YQ0sN7663ZbGXOYWTVUTYCGWnW1GxEHMfhw+8uFwHG8EqUzMzdw6PSNaG4lz85Sumrpsc49v1IpnuMw1VVRTEbzSmiY/g+RiZMrfd+vV4jovUG0Uhej314eDKSBCoODjBmvg1RSzIirPWkHMP7drHeI6LkB+6RSSbMmkBKshGJmC3pDPdkVoxeQXN5BUYEUN1MKUU158C9GckmICJmenhEJiCtNzHd3ffjuB5HJIf7PvYRc4vyewRkAAepMECSrLAyZU6byykMfhqnPlUmf4pw+e3bfP9EWN4YS/gmH7MjPtnD6xt+wj4/9ezC7/tDu8gbYbk8CdBfs2c8xXTGrjMeBgCoTFnzTYxdj8qt0V9yF1Ag5ccQwKAGtdO/PL80ROa8SrtpRgBSEpIpmQqq1IM89RpoapfW64jz9w7MoEIypnGGQpTnHZjrHCJUiEG7mZkCaGatKQARqOLu7v5y6d1sM2uqzGltDs7ifqJKz57JCI4jVK3P7jJAZgxkqLBmDAIVu8vd5XLZtr6VNlpUpdTP5d9ovR8jh0dEAkGBim2XZ733w/2j63F4DBHSXV2uqpcfD3//+PM/94fDv/Ph177f7V8sFovFYrH4m8wKoBeLxWKxWHze+K1/8g9FG6ka5s1VzQSi9uzSX9xvrd9XNqZCYUbM36wHYaatNa9MVqYVwM8Cr5AR4e69b6qaGft+jHHUr9QLZQzPCJLTNm06xjiOA5i13ihrRRUyxfrWmfBIjxSx3rfKr6fEQBRmRIV3SiBIqBBwjypa1yg2iLhnhXLauogex1Fd4sxK1KiqgHhkxJndkZztaejUBTCTLxUZYoAm0yN8eGWJOd0GmcnIDObwMRXUKhSJzBExwglJpmf6WZcOMoiAeHJ4umewrgEERkaSOUuwxBlEPuUWzn7fOPlTFZ7fQN6e0L79HF594isf8OVpzk9+3OE/yTHytm1nUvyWx/jkg1det/OS6l0nTU1f3YPMpPqsnLPG8c13rZynr6JVfdYzzc7ZFBaV0mKgmr5CnPXnsrxUQx55HlVmtRlGGCBClemTrpuuIgoxUYYjo4ryMieDinAuGiXnnM/6HYbWmpm0+i0AEVPdtm7lhFaYabMGpFTl3x0ZIohwd4egJgCWID1Yv0MgGdJbv1wu29aaqYIRI2OA0ZtuW996B+ERp5CkfqsgrVlZokGKauvtOnh4BtHv7s3MrHm6jzhICj3oIweuj8/w/Lh0v0i7/+p7733s22GxWCwWi8Xis8MKoBeLxWKxWHw++Z/+8S+nJiTBsWnPTbv13swpIrpt/e7uhanyeBjHnsdQwFRM5Xp9jHSd88c0gQqjxzgyIpOtNREleRzHGENEzKyZhVfQCm2mqip2S3RfBtBkuWpVtPcNkEx6EBBTgwiZmR4ZJNq2iTaIeDWeVSIzKg0HQGQERUTV/Rx5qEbgOAYJESWFiQiqShK1WSYBrZPKmstW7ot5uszy8UIAjUwfPsaoJDMqd44ouUb9qXgxpnNjjoyrIJsizgyQ1d0uo3QiAsMjSahWTj3Sk6gbNkUcOefXnXYOnLt9JYbmG56MJx6PySf/yPtk47dFu29s/NYA+pRXyHm7+VSI8bFWjSfa6ZfX9eT0nzgucEuWa6reqyFyyumRfvOMb58UEVPTNxLqVz5mBcvzNGSmvzCZqxQiZcTQBCizNn76l8/3zSl3BjMjZgR+k0DPp8Bq8UZ4m084BRhyqpwzkAFyVqrnTEA1NVU5TR8l0WmtW1MxkSbKTBXZtq2GFbZmpdw59j3dhRzHNX3UXE+SYlDT1ptIVt+7OtOA9dYrfjYVIJmBdGaowFTMDAAztRrSQMRIZm+NIBnkVG0cKWEXB6JMNyJQCfcRZIxr2tUvfXtkG96xRM+LxWKxWCw+T6wAerFYLBaLxeeZ3/on/9BEoWoQ/ejx+nd/rKeSRGukdsGz3pTMMRRkePp4+OiDiNG2y+Xusl0u2nrZnK/XK8jeu3sAsm2XiIhwkn3bLvd3N4FDorSw0vvWe+dZnT7zN+XMd7UsuLNjnZzmAsX1uB7HMGtmXcwero8Atsvl4fHxGKP3y2Xbmtl+3SMTKszZTYZoAiNCpPqeEoGIBEoJ7eEVfs30LjOPMR4eH5lJMDJJJPO6H5kAJILuMY5RpxzJOBPoitDUTE3FbIQfY4wRAqhqglBVs5Hp8/oywKSAWhGliELk8DHCfRqiJVHjFhljZEQyz9h9ps+3YYWJMkrPmYcFn/x5M2aVM8Sdkuv5FOJjq8evJ7pPA+g3hxZWM1c4hSW3DPo8nzd+9tbXP5N8JT2vuq6+uo2IdGmngRkCKGhyS4GBpyk2P8YqfWKq+mQk4Hm6rzxHRFtrtRQgJmIqZql1rYJMRCldIsP1fNUEVNBwG9zXK3GmRwXZ8ytCxWNEjNMCXsdOIqsTbZCutrV+6VsFvr23vvXL5WKmIlqFbVEIUgklwgNJNc1MkJfLhcAY4+GjBx/DFD6uPg6Al7t+d38RYWvWWlPTNsvUZmpmXdXMBAkyI4ZJJc0ZY4yx7/suQG+tt9aaWWvChKJ1y0x3J8N62+7u95TH4B55wBhIcQ+7e7BvfPkbP/O9n7H9mVM929e+8Y1PuluLxWKxWCwWn0FWAL1YLBaLxeJvBb/9K7/o93cC2OP1+nd/bPOkdkCYosxN9MWz++3uIiQ4kA6mmpmpmEn9Zr0HQBHJJIBmrfzKaq313rbu7hmZmfUTVkZNPLMxRkRJM1JEet9I5jRvqGmrWYjjGKXHMFOAyXSvwWfwcBHt2+V6vbqHlVYAwgyP9KjcWAhJwiP2/YCIaksyIt0DRGSOo/winNMQS36d6e5nBp6sknIkRFStCtSVuYOSkLkdKlUPNVMziHjEcHfPcjJEBlSs9SQDKLlzXU4mMqGis7ysSGB3z2QCURpoMjNZYwxjZtCZvJlHAKQgyJEVlQNTLow8B8OdIaq8qo5mqYxzZp2M7xNAv8KrDegptxBohdFnDZkCzmL2zWHxxt5m6fdJSA3MnvDLAxAK6hObc/1dLebzCKhEX28HfXoB52Feuw45A/QqYgPQMyI30ab2ytNE1IxMZiZYrzCfVK5r9N/5rppZdgXQKllrDjaL0qxn1/1Jqbg7SKqK1ledqak2MxEpbUi31qvirAK+rMKLaa2jREbQkSFkk7kUVFJ3ADVskzUvVCDCbtpMzaR161sds+rYta4yVwYiCELrEOHuw0RMtTVTgQoy85w6aKYKAYMB1kbarMQy+/DHEdkakyEIx2OO9l0ZX/Rj2//0+Z9+/etv3KLFYrFYLBaLzwsrgF4sFovFYvG3iIqhoYrLpVm/Hg/ivZkoZNta0353f/niixf97k7iSHdmEBSFqhhAZlmeUSVfEoS1rq2p6XEMH+7hpiYqVREmOcaITJARISJ96wAyOIYDomrNWiaPMY4xIlNNzFQgxzFGREQSUFVr2xgjPCpxy0xVieAxnEyIiLYa/Xe9XgFVa1GJeFRwyPCsSYkV9KlatWPlSa2YIIkZUaui8uJIQs/KsEBAYriPcUAUqP51RmREjSeUCCdErc3aMnn+QUT6CFWFSDDNmqjsY8wphWRZQQAkGRkZUxSSp5eYFZ0LEox8xXZR8XjeGtOnj+Nl+5gEtE6YuFmn8TRY5hlf35LppyluvhHyqijKKz6PlDeJCc4w9Bb2zp3Ml/qNNFtv4edpzyCrBy0vz5KomvUTc0VtpjOTlttlvBIjQ0rlDIFWFHs7swqORZBsot2a8FWTtQpBnD3nyDx79HoOKqx3VbvdJCDBFDK64E0AACAASURBVEkwhSmcJwmmqphqtcSTKSqm2tTay/qxNTOZNmdTkWpPo6Qe7ukeGWoqKplMRqSTIaQJSrgRmSXtGGNUwH13d99ag/Dusl0um5lWk741U4CRmQ7SzEBkpg8nIZA66ogZQFuzu0vfei+HOeX0ZYtADK2htYRE+PXYR0aCLsIUetqRP/m7v/9HP/9TD5eLPspvfvObr7+fFovFYrFYLD5frAB6sVgsFovF30Z++59+xWN81N7/w5/4P3/h//lluXTtQnQxvWvbO/d3P/aFF0gZ+8MYV0GaYjNjxr4/ZgQIa+38SUpFdOqS3X2M1luzpqr7cVyPfeqVn7gRzExEI9LdI7JZryLndT/OrjFY4/7mByGqvV/c3d2ZHOEeIVNhC5Kiam2roW/7foia9RYRAlhrGUGgWT+OcRyHVm279xFJwMygolq9VyFIlXJXM7Oi36RECjNFRVSjNBwR7vXHa2hb2auZiPQaeJgvr2UWusfw4zhm1xQ8K7PMRCT9Zb4pZM18I0moauvWemXKkUjUVXdRKetypc8CyeQRLgISEVmi4LpbFRVmcriXKaNGO543py6bpe/NafF+Ke84Q+3XXND1sJ0xZFZbuwq8WgP5XrV51Hw6IM7pf5VdykxZbzslqgZ+VqqlVB4iSoLMCnrllGbo+SggRFY7/OVZinbr07B8K/yqTq1zGaBHSNIIqRGWmCsuNSqwOsx1JUorT3rNBeT0nWMW8kUzIhjktKTMlBxUwWXbXrx4Xh3noF96v+vdrOb4SeW/7qGqgDLTx/AxmIzw4SPCmakKa81aM6sifqXoWdMF5ysjoirbZavLvbu737ZuatZMTZJ5XK/7vpsgI/wYx/4I8v7ufk6kJMs6LXMdJWe1GvHs7u7+/pJZQwvjGAOivd/1++dJfRjHHnRVMkFnZMixP/p/9Dt//OFPfVESL/7k/Xd/GN/KFovFYrFYLP7mswLoxWKxWCwWf3t59138+Hd/dvPnXzi+3C4NPpJ3umkztdaQpqq2dWXCd8tBP+K41vAxVb35apmYiVsyInpvrU/5xvXY93GI6LZtJDPDPbatm9kYPoa7x9Y3UQ2me5DSrJWiwHpn1TAzVHXbLvu+H8dxa/VWkF2hM0Ts9E2Pw9XMWssMETFrmQFIs7nDCNbgNo9MAKZlv2VVjplTl5E1VTAySWpSKrQFcIxRzepKnyPcPT2YpedIxsxgkZlZ/zzz3AjmGc5OC7CUibmm0dXLCRE5ZyPWEyHWrPUkSNyCYVHDPFvUlkSdQEBVqp0dmRGocPYWQEckqgR9jjdkPk2VZ3EbZas+w1cwMzHTYrnViDHj3xkGp0dkCJ5OInwlg+YcoDg/vg1OlNenC2JqQvBE5CGiYsB8rNrHZALQmk+oT1/aJx+Lmto89ROehXHUGgKBSIlUUpCiPNNtQigglCVP0bIui5SYO2+Vc1HgHFCoUsIYUWj9rRCgmW1b662JSro3la5qaiAjA0TONj1ARET4CA9tStLTyzPeZ/psAMy0tda3ZipgztssrGUOa9N0bdbIPPajcvpkhntEXHq3soP4IUTrzcRUVIjzlwFUVCg4l12Obdsul0swIJBmVE3qEZGJkULTIyMiEjiOvMf1q+9967/56Rd/P/njf/zRu3/p712LxWKxWCwWnyFWAL1YLBaLxWKB3/6nX0EGqZGyD3zhHQxvnhoEEZLZFd1MkTKu3dAUMi3FECCDEdGsi2iSfWutN1MNcozx0eODqj579iwzMyMieu+quu9HRGbysm0EDx+Aqratb5kk5e7+GQF3j0w13S6Xx4eHfT9ImJqZtdZK4+vuAKy1yPCI8FRVMyMTEBXNqQ2xZl3E9n2UD3dEBEFF65uqjOMY7uGRmMlzFBmiLaHH4ZEZmcdxRATAnHbrPI5xeFQrl5yl6RlARw0Y5Aw6IYTYrOCWzlqmmVoEWhbeim6r6svMHJGEiFqiLA4vJRsz4/Y4TdYzTxVRiEIwho9jABX5TjvwiEzGjNox+7uVm1beDJGcveJKdU1UEsxwiEl99ib3eGLTEKBiTVIrxifObvTLDHqKXGbmXmV3sK7/6ZvzNszw9lkRmNhNFV2BcomVbzGviJhpU0NV1gWiIhCCtwBaRSBSEzLDIxlCmKoE6a6AClVlWpqzvNk55ysmbF7EmeBXwq2q1gHJTG3We79sm5mqqZnqFIzMZYXWVEXSQzIlqUAN7gv3zLNQffpjAGx3m6gk08x671u/WDMRZaaqttYul61cGvUKSxXNkZkUhakQOPb9ww8/vHXDSzx9f9l6b6Y6je9kM2tqtfogotpUTMXkGKMq2K136z0F0JbgcYwRY0+hahDhke348M/fub8fTce/++73Pnjc3/v2hz/cb1yLxWKxWCwWnwlWAL1YLBaLxWLxkt/41a9cNnz52+//F//Lv/rn//iXj+0CUKi0REpXvnN/t3WTHH7sIjS1rW/p4fvo28XUKLCm2mzGqaS734ahmdm29Yg4jrHv1xmZNUvycDc1EQMlPBK4u7+HwN1L99z7doxjDM8EeI5KE6kEFoCJDB/uDsxycUQFeTdLMAAD1T1qCuL3PnrwSG3mNScRPC0fmZnVpw5mMPt2L9aPGoxIVgB9FplVVTzTI+b8OcoZD5/j6KS6ryaCTEawdAl6y2+zskbkDI8xhmdSVVlqjoiY7WpUQ7wE1qAQczweZ2W6jjx3BUHtFnPmXwXQ6dWwVUB02psFOoXOAlWIZMXHZ2JLwWklARNl0ZAKOXEKquudxPmJ84xuJg+dgmbwyRNK1YFaLZgfAbct6wWdBm4hBK1m5inUzFRNmmYiicBZZ06eQm/epCGZ7ke9e+pAIipQEpEh5Cz7EpIkE5iLCVWvnmc01RaomXsZqbWysfXCzCCSmdbUVE30pSIEBBHJyHD3KmqTFAqScXhG1HFVYKWUVmlN1cRMtrteywlaKzDWdWJShWUBI33EnGAZUW7o8CGC1u2ybabqHu5HZkzhtGpmfZFy611VIkJNTU1wTlZUQEGVkl9f7u/sckni4Xo87uPKBMTpoDgzH4Vf9HzUGHJcL1/7xjf+ir5fLRaLxWKxWHwmWAH0YrFYLBaLxesQ+J1/8LN//ndefPM//BLMtqaP7pWVNREVbcbLdt+3bipdNY/h+363XcwsAbEqy8r0Bs9GLkWkmptVOc2MajFPgwRZUwHH8PAkaVsva0cmRVB950zWIMGIuAmK59i65HEc7l7z/ea4tsiIUGmAuAepTEnPslg8XHePUFNPJjNIDw93ZBVzQUGZgLVtUPNgNUbDI5mJWzZ7ExHXj5cKsqLniHmWRE2hQyTDY47QywRBpnvVwW/S6WmMLjd0EhX7Jhm8Bbt1u26mjpld10Q9Ma0WrdhNwXze3duNrnZxWSFmSC8iU43B6XJ+GeJmyawz8mWgelOHTCNIiaLP16TE09MwUhvMbHmeOObsv6olAzLnGeLcW0XPT0vQU9wh036hs5vtieBpn85ZRJ/Z+0uzdcao/aiqiJ0u6Xodz6mJdZ9QETYqXy8HRUk06r/l1sBMis2a9tZaa3KrcAsFUJy35/SAk1LC9GSCLDGIivlwIU1BpAq62dbbtk2xhhpaN4LDh9jUT5ddvQrY9YZLD9+dlb4n6y2T6SIwk7vLxcx4vj6m2pqZ6XHsyRRBv2xqmqVPOe+NqomJmEKNphClYESMyAwO0D0GmJm2P/7f73zrp4+fvuQ97vI3v/7NH8p3pMVisVgsFovPNCuAXiwWi8Visfgk/sWvfWVk/uS3/uK/+l9/5zd/9SvAnirlN7izdn/3/HLZQOR+vb9sphoZEKjCTEvToUK9pYxStmgx0947eTaOSTGtuPZ63TNuXeAK7GYCeLlczGzfj6OGCR5HZgrQexeRMfw4dvcwM5FKHJEZ7m7aSBkjarBcOkXUrFXmS6Fao8AjPDwjlKICFYUpVCmVUJOQ1rdt24CpIq4dZLLGukVM28Qt0tyPY4yRQY/wiEhUJp7JDEYGI9PjGHtEBmeROQlrTURGVOdaqjtM0ZpkiFI/1FFuaWNVn+vaWit9c+utSr5PUdEaIxlgYObLZTLOWhAopcVUfDAyM8KTHuE+8NTT8WS3cobLYiqqgM4RdjOPfgWZagwkMMvKmM++baygIM+zn5MPSUYkM5J1QykERqJe/LqWM+CvxnSJJQDq2au+NaDdq2lutYYwQ+FTVlJnoqram5VEo5k1M2tqak1bN1MFkDEqnc5wAUw00sEQQE6NdzCTqWIEPGKMUcswvV962wA0095bxhCimV4ul8tl65uJgEhVJDLCRQ0itVozjjHG8IhMNlEGfXcVVRNVU4VOEQtBVj4eMbbWm1kyzMxMxzgIiGnfuppBplU8CKhZ22DCTAfHOAZzUMUsRRAJRjx+9DPvfetPf/GnvvtFH9i/e/nw61//y37nWSwWi8VisfjcsALoxWKxWCwWi+8PgX/9n/zcX/zY3b/7uS8JWthuYmJdoRU2Xnq/v7uTiBiHIAzszTJG+DBFCZvLbFs7vCWSnJLgqu4qIJmIYLVsa4Dc48OjCJ49e0ZgjPHw8NCs9d734wj3jDRrSR77gVMjbWYiEhEArLWsoq5qJjMynSJiapEhoq23ahunIDPB7LMYqoAk6LPmKx6J0vyqEoycoXImASE5Dq/P+IjhU8ucmWOcmXPW/EM7jhERc/ZdpkckUTFhBb6tNzUj4Zml7IAYoIHkbLxSRbZ2KUnEaRjWam3PTFm09w4ig2UhYbIEEcMHAaqk1CxCMiulRE6/91RXo7wZ5UJOZsSpCXk53a9+rHb3JFV11q4ps/x93vPqAc+MfXpZkLjZMl5uWu8TBYXJjLMELZVTi1ipt2saIZO99aaGxJkdi6qoPXFUn6rsjGAGWA+JqIoKIE21mbbWKpM1MwHI6XNRszHGMY5jjIr1e2tmCpllddQ+QZuabZiJalXxA8zWupmpaeTLeF9FWmsQEcW29b5tW99yKjSIWWAOVVHTs0A9XSsiUpX/NvUbYqogY3irmYGZIlCTrTdRkGkiohCgt2ZmUQ4ZUxWJiMPdto4521Mg6rAj+DCOKvRTgQCFIhmSR8oF+3d++ve/9HtffPZH+c63P3z3R/HdaLFYLBaLxeIzRvvrPoHFYrFYLBaLzwAC4F9/E8Bv/OpXUhyQQx9BsRAhXG0/4mE/tt6b9aZbpsfwdA8fAqqKmUY4MudMt8yIqPiyAugkzbpZE2kZjCQBhYqoh5cqYRoqIqVp61v5cskQU6O0LmXjtWYVQLuHyBlAA2Y2I708pcaEitTnqzwcERHexJqpqdURPTOITAiQSaYTSmYMj5s7o0wHw2NkRI7D68HKTKtXDFJJ07a1Rqdk1nQ/gZFtqiBEKtpuraspiBERSVETNYjmNDpIjezr1gAkU2cy3oJZAxQr41RJJilU0XoEIpnhvic5HSNzqqFN33LdkOlRhojJzJRRBgyeFo0ZLgtmH1oRSUEiiXJYnKDkFvnyf2A1jc+wfAbQFJSEYy5RVAl6HrPUKhBFlrSjVVpKbltv1gCZITqoqtb05sQGyYwYAjOANZZQRc1UTAUoH0XFytOpMvP6eamZ1KAZAAoCRKaAzAxmYsbQmSolqLbWrGwioiLaW+u9t9ZKMi6AmfZmrXcykmHdzESVKpqZY+Tw8OEjQlXVbLbwQTAFUBVGCtF7q7hcQGSaWG9mJaYRisi2maiQ9esIqMwZIpJgVdTNtDW1Lr1rb9CWicP9Yb8eyYMEEJFCagIHgHe++t57//U/+Okv/WQ8+/CL3/mF97/2r35E34sWi8VisVgsPnOsBvRisVgsFovFD8yv/9ovAV2oR//ed778O1/+43/UhxqMMJLG7KrdxBSK8DjSR/roJs3ETJh09/36KCKVx0UmRO7un239TrRxBpgziLxeDxG5v7+/XC4i8vj4uG1b7/3x4eEYIzO3bWvWVFv1bVNmlMlkRLh7yROmMFjV1ACQbK0zMY5j23rl1Nfr9fHxMSMFFFGW6IG5H34cJcyIzIRIToXCkz4vWIqPEvJWqBojSOl9IxikVHl22/brNTxUX1Zu3WO4azNRSaKpVom7LBxtu6g1UeOTCYRMxvDSUrh76RK8Ri8CyRzh+34wUgFTS8/juosIgSBHjiN8hOcs1LZyVOSto1sab2kiApXbBMMqWwOoGjIqyDXznIXwGckLZqp81p15The8CTmIc1hiiUCkpMNSs/VUpJt2s2pg6+mVjsiaQ9l7V7WbP9pUS1IdMQCoadbpMJupAuHerN1t2+WyVW5LVk24dCAEERFjjCoX8+ywRw4Colq+l9PUTZO614mMqUGJ6L0/u392d+nNNInWTLWBMLVurVQrALfWeu+9t0REHvtx1KKFWcvEcYwxIoKiVq+VqkBIRq2OtGaVs9/f36lKZvhxZATIbWuXy3Z3d0cwM24WjrPILpkZkSNJUagRgtak35O5u1/3x0FxGIlE+EiJ6/s68Pf+4MWf/L3+8IV/+90P//zR3/v2t3+k33cWi8VisVgsPpusAHqxWCwWi8Xi359338Xz7/39Pp7dP/5EGJuD0UygSVLMcNet90tTmKTE3jTuL83MALg7CFQtlxmkmak2lelN4GzbIiMh0swq+9v3Q1XMLM7usZy1V5kNWEBmkgiIqpL0iGMfgIiqimSmezZrmdz3fZohosYA5vABQqfFmpExgj6T30oZy+iQZqqiBJlJwKwJ9JyzJwAiCWjvWw2Dq+PXyYM0tbMCnO7h4WImIgLNiIzISPcg0LcLRcrUMTPukjX7aWiefzMyADGz63Hdx5GnfMKsSSIjVRWCyBwMZ6k/FGIiNl/w25Q6gGdUXK+qAEqUDBlARo0kJKfOQlRUVTKSmVWUrhGEckueZW5WOfjLBvRLAcdMocsR3axdLr1cLdPgMd3gNdqwTk8yPJnnD/eVYmupNAAJDy1TiEi5SkTw0v4yR0ay1N2ZEe6ZAaCpncMXw0xPPYeaae9VcK67x8zUMnjcxhRKLQxEa021ZVCgqpZVRI9AheiqRCS8JjkmIUBEjmOYqKpBVbTWTmgKtRJYC0AmVdD7JTJ8jLu7S7OGZO22tRYREYNghewixBR3q6gRmqoUG+SgPIyRzDJpR4YjGXb4oZeDh4zLh2M78IUPvva1H9X3l8VisVgsFovPBSuAXiwWi8Visfgh8D/8d/9IE0ixhDIpCbQ5ji5la3x2t93fXS53/a5xa62b1hNrvByZ5WsGAIiqiCgFTJQJt7LGCj0jKrmeI+xYJU+PcQwRqEjlpADGcIj01iNi34/vffRIQkSFiMzwFNFMHmOM4/DhGdGsmenImOdBZqRHpCjVRKy6uzlH/nEr+4FIZJDc+iaq5IzBS5dLqKpG8JwnWPYPCqRpFZ9HeNSEuiQhaqLHdY/DS+pAYrtcPPI69pw5uEy3RBBRkg3xiHE4BaLaW394fNjHrq0l0zNFzKQCcyHhESlJAcVETa1BlJCSUCcy59S/m0VjxtEK0Sk3RllRos4gubXeWlNTRpZl4rXxg2XqqPsrIjcFx6nNOJvQwPRhA621u7stIzMKz4zkvMWlzlbRCM90zhusNlUsrfdOYt93MlVrJKMkM9zdh/sghGcQPoUiTCCrKd9bUySEgmzNttakXsdm9/eX1ozzRQIpVsdrjaC7x4gxYoyhqioWzqzLFMmku4eXDgaQpNJU9Ez2mZkel7713iEQhRqa0gxzhQKIiIwAYdbdfYzx4vmL3jtjLjmIoLzXkSmmrbda00mx1jfb7ikyjvFw3R/dh4pDUoDMFLgf/eGLcbmGDiKkxW9+/Zt/Zd8/FovFYrFYLD7PrAB6sVgsFovF4ofJ//jf/ucELS7PH7700fM/PXg0CpqIqDa5qNzf3d1ftru77VIGBBVGkAHG1pqKRLiaqlqJAjzCRzApRE3tUzsjzfmjnCgwhj88fDSlEWeMeRxjuHumio7D3//gQ0BULCJEVK1VqioC5Oz6zm5uK4uvoiJPD23d+tb7Zq2V5+HMEiEqzbT601pT4DIjpqsDajUgcQz3yAgnRNVqJKNCIsIjxjHM1Jpd9z1JM9s/usYI01aF69a6R+7jYCJnUAsm0qOb9dahWv1lMTUzs7aP3SNabxRJcHia2v3l4hHhPtxFVVqppYUCsS6iSZZfIit9FjCZZW0GBWJiyWBSABMR1Sp3k9lbU8DDS/+sNQlwCk/SPc5K9BwzmNWOrnUI3gYFMmPKPTLDzHrfZmc4nZWoRtrZiG+t9d7LaVzvhyqqq5pZz8R+vX7wwQfJUJVt62Ugrxl/dS6q1lpX0WrNq0pvrVmrkL2ZmEpTsabN1FTJiPB+6a2Zag2sbGYtIt0DOkdrHvs4DnevtwJB8eFjDLVWOuxqY5tJDVtkhoiYWd/a1qxrK5u5qpJJRjOqkMhz9iPGMSJi61uV+o99uHtGlApGVNtl61tLETFtbSMjkocHtI9MFxlApKR7AAeHH6bPrh/9xDeff+fn7PG5jbuvvvfej/qbyGKxWCwWi8XnixVALxaLxWKxWPzw+e1f+ZWjf+Q6iA+e7x9+9Pw50HCxpqaoYXm9X/r95fl2d2/KPB51XLvCBGBUAxbntDv3cPcYrqIQJL16nTWPrpwCEXHs+7Qo1EOU6z4iWTlfeH7v4bG1vm2btVbS4LORKwLVKZZQUYFOBXHloOGhampWXggRjHFERnWvAbSmFYuWctrdp7vDEyKReb1es6zFoqWpOI4jI1T0HMpHFQVw3XeCrTU/PD0FkskETVuJm8uFMc+dkpmmZqpRQxJFapJdTXck2HonEMwxQkUv21Zdb5JqWheVpGdShIIyNhMQ07In14t6lmq1Wz+qO5wwM2vNo4wYwDleEkyAbbbFqaJkepXcX5acWbksWW4MNZNpu4jSVBCgmV7axvOZcs4/VFOz6iNb6w0VmnOOAyz7ioiSMsZ4eHgAaIbW1QQizMx6bk2h7H3rrauqDyegIr1vCs1MVTHVZgaQnGMHk9m2BsExjmZmramaux/HoExNy3Av/XeVrZPMCGb21psqBFY3wCBmaprMMof06uHLFJVk0sdwH62pCqZ8BICgLDS1XCKCcRzpwSRExdp2uRMzmKKZtksSD4+P+9iHB6yhtQQZ6cB1RLt+GP1ZGMbd93i5jud/sVQbi8VisVgsFj8UVgC9WCwWi8Vi8VfIb//KLx69p1ps2/7soz/60u/+/P/7X9qLCCibJIyQzfTSrKVvSM1hwvThHkyqmqkl04+xP14vl4uq7Md1+BHpIgqRpNwSOQUUlHRQAb0Op2jfLqpG4hh+uVzun93fPbsHEBHWrGJfQEW0WyV5GjWYbsoQyMgavhfhJSJ+vD64DzLdnaziMzLjer3uxzGGmykI9wQYkfuxq2prvfeLNSuTdWTUZoBU0zki9uMAuLUOKEl3zyRBFRObddnpsRYVmb7pzBxjT1DrEoAyMFRKSzCC4QGimYU7ydP3oALxqEQ5Ys5SJERb75WnqxiBsj2LaO+X637sx5FBbc1aOzxIMdXho1rqRArYTDP+//bu5dfW7LoK+JhzrvV9+5y6VWWXXYUdmWDiAJIloJFGZNGgWqBI0KwOvXRoIFki/8H9C2gkEg136NCyO0hEREJIqR4dDCIiESAnJCR24vhRrvs4Z39rzQeN9e3rKEJCFpbLj/FTlVS3qu557H3O1dHYQ2PGdLd1UDHzjJ5vmx4ZsZJrXW+oNwBRtRJ8AKrSzfbWZV0lVNEV2jZbRw0LIgJVWbm/R3isAer1d5k2QCJSFWYwjd60mUSEiLTeTcTMtr7tl721NodP94jobRfR8ESViDZr69GI8EKpauttxnz2/Nl6zCGyXnwouY2EA633J0/eyEyfnuUKMdG9W1fVdflQVRRmTa39xRdEqioiVBRVx3Vcr9cxRu+7qtb5CkFVJQCgVKBaahAVgShErPX98uTNN6/HeBzXyLqO6YUjM1BSBcEUfbJtT/7973z37/z89UnPCPXxpa9+40f+hwQRERHRTzkG0EREREQ/Ik+f4uPf/dyW91Z/8xtv/+3PfPgfbZaoZmpWlPuGutv73noTiXF9fPmyIkSgqMrwMXozayZApEdF6121iWhEquhl26tKKjfVKkRBbFPr2lpr7RaAiqhYM9F16g6Z6TPmmJnZ21pR8MhzeSPCKxMFFagAWatcPMbVX4WtVRlxu21Yc845p5mamaq11gCMOUWkmVnbIFKVWBsKAFaxNs+55DHGrZzbUOLh633c7vap3CYmck1Bq60LeB6uZtu2reKzQM755kwRVWjminT1PFoYqbesMzM9M6o8YoafPWOVzMqI8HVrcJ3HU4h6pGethxOK4SmivfXjONa8CSSBMpVViF73AFtr8mqD47wTeN70U9F1rXD9wzoaGZVbs6ZqkDpXt9cncZZ/V0693o7Hyp5j/bo1A6Sqeu+qBmhr2poIXKUU9er39r52q621piJz5nGMcRxqvbLGMSLWcvdqS0tmiKo2c5/D55ijzk9GTNVUISVSKqjzdKBd9svlsm+9r5Oa62WS8wtQRATff3jrXMSe06/X693dXTN7+fLh8fFxHHPf7sza+jKAigjWM9O6WbO2mbXWWjO1jAzAI66RjkJJoDJjFgoxYn0H1OVbz7fHuf3+N59+FH8gEBEREf2MYABNRERE9KP29OnTN65/3P3B8tt//sb8a3+OyCYRJaKFNXdwt+3INJVNS3JWesUUlKmY2TrCZ62pqEIiS6HNmgAoqEgBVQI10abWXqWXa804M1VVm1ZVuI9jzjkrs7V+jHFcjxVMz+lrYUNFTCACETRrrdn0mZGZuVLO6fMcXjbzcJ++ton3fWuti4jPiVuJt0rOHQ05x0MiIuK8ejfmzEqBqFoBHr6OEKqKrOUNaNYtfs201lW0Ch4OQLVFeBZU9EyW3QVqYuuO4MqkV2YNAWrNiVSJeKZHjDlXpQPlqwAAHthJREFUdg7BOsC4dh4gWEluZGYha40nm5jNyCqY2TnhXFUokdK1kQ1ZYxfWm5w/f68cWs26rYS51sizqwggmeeEtpmaQG+XEOO8/QgBIiM8VmvYtK1idWaKiqq23lUEIq01Va2ENTMTICqjMtcyc1WqmtwS8CpE5BjzOEZrvbLmPJ/oiFSVlUGLiagMH5m5jmGuwZZ+XimstR8OMYhmYd8vl/2y9SYAMioTleeZSgiA6XPMWYVKVFa9CqDv73prD48vfXoWum6qJiJiqiJQmRmFavvWtq1dNqhG5BjXCA9RVHlVFuA+Re4D9/3TH9R3B0aVqMq/fP/3Ppo/AoiIiIh+ljCAJiIiIvrIPH367psv0abcP0K1XrscL673mRA0RV5a+9j9/s4nP7btO3JIzvBZGaJiZtqsMqVKCiKakeMYpk1EjxmiqtquxzWr1PrDw8sxjopYG8VjjFV9XfnscRyrYtza9vDw8Pj4eNl3FYnMFbF2s7PWqtJ779sWkag1mKCZ5e6quq7h1W1BorV2d3cxNQARAWDtMq9t4jEGADM7jmMcxznlbObu6/+s1c52X9nr2ZUFRKwK68POzG27bH1XtTGOOeac4R6ZULVbAJ3Ite58xtaJWmlyVs3wh4eXWRC1GTkzPGKVgs3E3ac7kK9u/a03suq6rbXtctn2i3t5hkdcLhdRGWOsqFshrbW+tdt5wL84wAGUqnaBocR9+BxzjrUncj2uQJkgMgTrmCHOS4krx79dMpS1x7EOAaq+eqDOfWfVFYvPOV89gKvlnZnh6R4ekZUrWI8snJvjue+7qkaESmXE9Xpkugj2vUMQ5YVUs/1yuex9601Em1k3VYUKVCFiqk3EULpeqFg179t5yrPsXFVjjDFHpZwZdCEiI6L3Zk2mH621bdsqgLW6oYAggTKR1koVIiP8GummAkiWwaFmR973Tz+v72QcXe46WrfXn77//o/2G52IiIjoZxoDaCIiIqIfC1/+tS8M79fCsz7fnE8wXU0vvTdrm+nlbt9620ya3kqsq0MaUXNGzPTISEAAzRX0FabPOdc08MyMjFgzCmfirOvwnbW2rTmJ1vpaFlactVZRExVBZQWQqtJ6730LX4GyRqyx4rOerLrGomvlyK3ZWSJ2X8sT4Q4AUHdfRewVE0fEmrdYqXfv3c9zht8PoCNiTm+trY7w9XqNCNXeWze1OWd4ViLOGjJW0i0i85jzmNa6iGTlmnHIKqhk1eP1Uc+Dda3WUcS1TdFaVWal6vloAK9+fBbIutZogByHe0ahtm1T1em+zkeuRrOZrq0SWUPS57jJWjC2KqlEVValnE8KMlNXfNus3XZXbp+NAKhMVbXWAGRWuFeWivTe1scZEeGxZpQza4xj5dVi6hHuLrr2UqIqCyKiHpmVzdrqO++X3dSySlHrK+CsNpuKohTNrPfWeru7u/TW5hioXM8/kKgCkFHHET4jbl8oEFlh9K2RXzhXRFREzhlznDl7VmZGwa211raI9dKBWVOoRtVMH9NDFapZEYLITEXPemjjS//hD/7J3/3Fv/7GmwydiYiIiD5CDKCJiIiIfoz8i1/7wh6bJTT71fp9Hr3UtNb08a62denbnfYOEUNiXmseOa7pnmc+JyLtnEhGhcec4wz9sszMxNxnZgElar1vl8s9AEDM2tokrox1EA6i6wwhaiWVadbMWkRUFiDuWYW1EpFZVSmACKZ7ZQKIXFvScVsAWQ1o8bXtDJzLwpGoQpVHqGrbthXUTvczqVVz9zGnqYkgK316ZALatJloZFRBIJFrduGcGFa1OeY4Zm9d1CDobRMVj1jL1tPdrO373veLmEVWRADVra+w18xEBFK+bgaKCLSALGRVRB3HiMwSWSvPkWlSqBzjiioVWSMeK3LNc6cDKIEYSl7tkdir84prVmMtRDfTprhtd6z9EAhUVdVWdj/nDA9UtdZXAO0+55hzDhHLLJ9z5bxishJ2Na2s6aEiaqZq64PsvYuKAH3bzkr1LQ7WtcK9cnDT3vt6PWO/7GZ6fXyoDFRB1mRHoCo8rtc5xlwvSOBsYcs6OInC2iRpzaw1FRFRWJMqNW37XlWRWZJqZtq8NMWGe7j7nCFVgAs8gXDvTSx1cxyWqK/9+bNvPxxf/YMPPorvYyIiIiL6PgbQRERERD+Ofv2Lv9LLrfDzX//OP/w3//lL//SXenttM0WZK7xKqvbe9iYXlU0L8xjXhyZqt+3jqtr33kwFZa2r2rrLB4hpuxVQRVStbWZ9bWWcZWTBqhuHr30GmCiqrsc1M9cZwIhcYxeZtW7I3RYzUgSr2jznXBvE7j59esS6miiCtb6QVaKioiqCQmWOMaJSVdUMwJhzlbW3vkEQkXWrN69EFDh/+y3bRMZazLC19IyCwM7sVFXEVLRQ071E1NTMICjItu8QdXdUCcS0rWa3mQHlEWP69PCMiMwojzUlXREZhQQgUiipVCRyXB9fZoaKQiUj5pjW1p281lpvrfe+rQ1owepMo0RKRCDWmqodx+ERJTiXqzOPcaTn5e4OgM8V0JeopGd4zvCVD6/n8byIuCan1+ONMJPWrFmrzDnnvvVt6733iMhIa7ptfb9sa+Ujq5BArcy9gFpnEVXbGtQOT1Ep1JjH6siXIiLGPNaRyfVlkJHrczez8JhzjuNovffe926ZtZrvaqJqUSHW9rtL3y8iNvxIz0w8jPn8GC+PXAcpK1xcgPHoB/DpdvcolxAtsfyN3/raR/WdS0RERER/CQNoIiIioh9rBXz1lz79vbee/O9ffMesZ0MbiK6CjCwpSEUDumSH7vu29623bioqJRWCFLn1bVEqKoDPGR4RKaIJ8aw5PCJVbeWWqpqZPj1zpY+y9U1Vxzgysgqrvyyia7E346wzr5kKAGZWVXP6tm2mOtxvhwdVzVpr4QlAzFbBWVVX4Tlv9d41uDx8rnfUe1/9aKAAqIiqqapApdYDVcC5sLwScFGgKjzXPDVW3bZuVwBFPCIyRM5FCGsWmcf1WD8iV6ISmTWnr8i7Ch5xHXNNnazYugrTY90khKqoKKobTCrmUZUium1bawbIGmVeVDRv8yOvBirWecOqKkhWXa/HmB4VrTUVjYw5PSPWace1vg2g9ZZZKNyGLACsFwbyNhktt3GUaSq9WWtNRYBav9y2LTMzQwpmYna+AFCZc3p4AurTPXzrm6ihZKXw4akmK4MWhZoUymOOOQo4V1lERKTOZ01vz1KuB6O1Vmvbee29mOZ6YEVXuD9jSkpUTY/Dc2aiqo7x6Ll/2Ov1CLMoBV7/0le/+iP5piQiIiKiHwADaCIiIqKfGP/qn7+rgVrxqeZF57MhLTIrBTCRTaSr7tt2udvvLvfQpiqi8ONIn5XVFJr5+PDcp2cUAM86Zj5/8eI4RrOWlZnZe0NJelSt/rDu+26t+RxZQMGnQ6T3LueCxEqfZds6gKrqrQNwz9abqnquJWWtKrPWtx4zC2htvccSkTnnnPNVPGutA5g+s2qd1MvM8FgTEPqq91xSufrcKwSvqvPgoZoIZE5XbWat6rxxl5UQMbMxxhhjrZVUFZDT5/V6VRGBRGR4+vSHx2tVmZmpZtYx3ayZdW0qYgWZ0xMQXcGtmmBr1k1WWVsE93f3276bGc428hkGrw9gjjE9IhNArg+yyjPdfQyfc3rG5XIxs4g11FyFMjXV5u4i0reOKlXdtn21y2/j2qU3IhCBVKjAFL2322cUKtj6tsLwiojIqlxzIpk5xnSPKqwrj9u2qWglIiujKkpN1ERVrZmaAuk5h89CQaFrXsOsziI2VGBqrbUSAUTMAhqiBXGfPseYI2s9ST0BidXVTvP4zsPDB7/wjU9+5zP2sNVjpaMd9htfY9+ZiIiI6McXA2giIiKin0hf/rUvHIFK1OO8e/YwPvW6KhAqiqqtVKSQKQooMisMsvXeRTR9Xh+6arP27MMPhru2y8NxHMNRlZUi8vprr6lqzLg1oNFbE5UxjtVNtrM/C1tzDK2pqprqrU2877tZE5zTzNpsbR/LraArUBQiY/VzIyvDM2vbttaama4KsEdUVlbJuraXaboWmWUtbLivuZEV9lZVjWNkZe99TYMU4IGZVbeoujIjwqePOdzdzlVjyfTIiJjNmpmp6RxzzinnAkaqqJlpb73vvW2tWUEq14yzQKREV7i82tEZGR6RcXe5A3AcR5wyM1b9eS0sZ2ZkhkfrrbWupmuQJLMSCVTvTVTWScb1EoRZa9YLEIHZeQRy1aKrqvcuwPmAn+skMJVuTZCVIYIC1mN4ewQrs3z6Ol+4jlCulB+FFUuj1uKJma7TjKKilRHpGdl661trplk5fGoTaSJmJVVq/XJvapWVGchSRWR61OOYHzwcz0cWbOtmIrLuMcLE5pDdxtjvX8MvffXlf/r0hy/nox3Xjz//ylc+wm8+IiIiIvoBMIAmIiIi+sn25fc+H0+2alqXLhCpZtlCZ0wt8wpFZQGZaeskX2Lr7bLfbdYeH5/PMUstIrNKUBFRwBuvvdZUI9Yacq2sEajpw5ptfVv12MpaEeWrlq2ZRZxBqpkBMt0j0to6l5cZAUDODjDWvAYA9wDOH05vG9byaqHi+4f7IKZagqyaPsM9E2u8AiUFAeoYo7JaaytsjoRnzdvFO7m9A/eI8MpqZgBQeY5IqIhIa+1yuaz3vprUq7675iRa31rrInBP97BmJfDM9cuIFAgSY3jGio+3rLxej7Oife5trI9bzkXszMxs1lpvrRkKqBQ1VVFbCxZnyA5g/WtVa61BEOG3H+tlrYCYWVZFeJ2he6FKIb01BSpXNu5jDlXLrDmHiIoqStZHsma4VRUrXT8/dahoVkbEmoJem86ZXhBr2noXldZ621oponJkQEX61rZLVo7H63GMVVfPyIkKj4eRh0elmJiqRMzd56X9wuzfSzlEm731oT2Z+Lk/ffr0R/RtRUREREQ/LAygiYiIiH6qfPmfvZsSlQisZYncu77zyf6tbzw/2lYjQlQLkmIVilK1srbvd9v9/bZfIiLmeHJ/WfsLIqWKblK1+sdhZqtdW1XI788uV0FEem/ucRxTTQpYI8WegVJUZeY4DlnLG5EomGoVMivCV5L9+Hi9HtcxDkBRyKqMcA93F4GZqepqRh/H1cNlHSMUE1ERhcLdK2ul4gCmR5TkOdmhK2HWWylYAFNb78TMWm9975lppk+ePDFrayF67UtUVXiMMc1MRSLjeoxjzG3rWTXmvF6P4xhzuEKl5Pp4ADAzUS1URIr8xRloxW2p+QyIZR1K1N56VVbGGo/Wph6zMkV1BdC9tarKqrvLpYDr4yOyAIjKvu2996pyn3OOWFFzRkWi0KwpVFDT55jjer1u+16Q6/Xaetu2vbcNQBX61tUUgIcDtW3buh6pqsPn4+ODqZmamWVFAeuAoIikyuX+ycfeeuvxuL58ePH84UVGRGWoFrREKzIzMWNK+NXvPPH2Pb71Dt59/+V//Ux8714zWl0aWtOPP33//Y/se4mIiIiIfhgYQBMRERH9lPvtp+++fH6MwHeivv6Jy9/4ph/XA1AgGyRKUgXazh1ftX27fOKN1/emJoV0lAsSFZnhPs2stzbGmHPGdLMGwN0jo7JEzqZz690zHh4f147Dmnd41cNV1Yq1j3z+OBpxhtnTPdwj4kw3zyZvzDkFaGbrnF4hI7PW+HVr1qxqnTjUyFhbGq2Zqs5wUVProrp+m5n21i7bvoYvBDgnOAoQVbMSQKBi1pqoHseY7pEB0RWpr0Z2Rowxp8dKuguoSlRV1qZt07bGjq1pYdWL7RhHZu77vpL0NSrtPo9jVGa31loza621iAiP3htQEZ61/oWrmqmpmU+fc/ZtQ9UYo7Kq1tE/UxH36THCp8cUxbb1iqyEiSkUJdBajXUxzcpjjtbOU41VlYnW20rVC6kqfdvWkPQ52CGi1rdtv3/tdTOdc37w4YcjIk0LGnp2uiPDM6WyBFUZIiY6vfzlw53/vG/frnpQU6t7vP0SLfDZP2THmYiIiOinDANoIiIiop8VT5+++9aLbCPuX0ZmtLhcHj/17I0/AY4MK+3apaBWcrf1TdFUmpmqabPeOxTpYU2a2Xy8juOY42jWADnGXIFsTI8MFPq2RcTLx4femqnl6ucKujWpFdQCqEwUqlYgurYxzo2KbG0Fy7aC3fAAYKprDQLAGqe+9ZmRZ/yq56zxGUDLCm3V7Dbwgaw01cu+R2S4Z+YasvbM6TndtTVVrYKaidr1us7vTYhWISs9IjwyogBAKtcsxvqA1UQ36Ka2NTNTUY1KiKjp4/Xq7r13U1MVABkZ4T69Kk3MrKmaiERGRopIVbpPAJk5bkcaVS3c55y993PnxGPdcrxl+pnlGe4x1PTubs+ojESKlApETMz0zO6lRoY1W2XwKimoqpacKygiYr0BKFRUipm1XWxbCy0Zfozrs+cPMyNUoAqzSJgIKhUeri9H+6M3f+evxWfv6knOwNjg2vNNFpyJiIiIfuoxgCYiIiL6GfXl99479mehx2wvqwC1T3/zxT/6zf/2lfc+//jOE82u0pBwVFZqE5OSkm669aYFFMKrb5uIzZlAReT18SF8aua27xD4GNbURKuqNW297a1V5hzDVAFEYs4ZlVu/rMTzlp+W2XnTUNb48E3diIiqtGbTx5wDqmtPeU1Bi8o6VzjnLJSIuLupbdv28uHlnHO1jN09IkTUtM3Ih8frh8+eb/u+bZu1LqoCcY/p4eGZgAhUcnWnK/f9ctnvjmMA1Xrft23fts1MIjWyKVax2sOjMirHnD69qtbS9DGOzADQzQQSESjJQoSfu83n9nWZmQjcYx0tPBvfqG3bRWTOmGNmnv+bqtzdX1SRNSNTFNu2VZZ7zMMr1mnBStT0uNzv1tqsUlMzRZWIifaCbNv22pPXhseYM9KP4zrH8ErPzJQAoBtEkBE+r+Mao+33z77j9594sq1JDXzts3h274EP9fkjxoeXb/J4IBEREdHPGgbQRERERHQq4Hc///YH77z2R5/7hO2vvWmvvcCLRBTKUsqkREylUpAVQIYgK1IiSgoikIqt6da31+/v997NBBnIyAyREkVXQ2X6zMqqipI1XWzWC4isLGQVMk2gt65zoVaqDJF15S/WYrKKSEVEpAMSEXO4iKioteZzZmZrHYLMHGOsE4h1O8y33nZlFVClMIvIMaaqmJo1Wzshd/tuZgIcY3hErfFokVVGFrE5PSNf3ekTSA5PDxUFkJXTfQ2UZGZVAqKmIjV9VKWZbr2vrPy8tli5lqIBZMEz9m0z08pade+CFAq1LihKrAOPmVXVWtua9a2JAkBmQmCtZ2RUZcCst7713jzjen3ce4diDF8Pt1dFYM70KC+UwCsrS1UFVRWZBalSUaBg8EgfeNxyy9QxAd0Af31/6wUnNYiIiIgIDKCJiIiI6P/q333xVwZGICYG1r6yCFQAEaCZfPwN/cY3PUe4ZLiIAplmooXNcOntbtvv7va+35k1EctKlTQVxKwYEV6Js8aslpCIikhfR/kym5QCVciqyoyCqInacRxzumes7Y2qWHlyVvqMcUxAVLW1fhxHROyXi4hE5DiO6cM99n1T1TldRdQUkMyKQuubqGTWql2bSkyviDeevLZvW1N9uD7OOfNcitbWWhUiMmOdaIzMzKhKrJRc0VaJeYYXoGbrVqOZ4TxAGKJYm9QQhEdmrr72ObVhLatm+ta6qeaqTqvEulsIqMhtumSl6mnWejM9n6y1byIiWmsExZq1rW1bV53j+vz5MylP9+twIAKIzGvCAxGaIqPSxKRg3SzQMV/E/bPv9J/7x199+hS/+vc++9m37moUouD29P3f+2i/aImIiIjoxxADaCIiIiL6gf3203efv8g58uVjRJT4fv/4zp996r98KrZrfszGsNZEpdQyq7Cu0KWhukErmpqqNO2lUGsQPB6RiRTDbXFjbyqFMWdEZiVEet+abQ+PD9fHxzmOpmuiI4GsyjknCgLNtZSxCsBAolZTesy5GtD393em+ngcpmpmIrrSW20tq3x6b2qqlZnuiLhsrZkqcMwZEVGpqmJWlVkZkQJ7tUxdCZQCKmKqBkihPELN9n338ETtffecnt63rqYQZMQKndfMSGttzYy0bVsXAlGSWXPOtXx961oLqkoAkSgkcH5UUT5nuFdFRBUqPMMDVVCBasJMOxSVpemFqswCyjIELfLBNvi1pgHYc3tR7cmb7o+ZLsfV8IkX/+PPPnzRP+CAMxERERH9PzGAJiIiIqL/X19+770XT/602YjtcfOO6qHze9uzTx5vRlRVK4SoqKQVStNKRBQqalIlUTK8sjREpaREtHTftOmWQK3dZZXeW9N2HMf0KRlSJZmqJRnrUl9VvTpQuKrVgHjF+mVkrJJw711V3B1Ya8gCQYlkQSCq1kykKiMyApWtqakIEJmR6RmmqqaZsU4mvgqf11YISlW7aFexrIqIrBIVM/OMAlrrWRmVomujAwLoqlRnAbDWItzdW9tS5eop0HP/ImN9AKsprqJQ8ahrxhwjkT5neFSEVEFSsqCKLKkqFSlVlQCaiHhCkK6oF2/p5bu//DX52mfkxSVEMssTiNK0LLOmqbJd8ulX2HEmIiIioh8MA2giIiIi+uH79S/+4r3vmtp9q0JBREqlREoBAf7Kn7589zf/5/tP3/36dx4tskpHGgpRklVZ0kwBiTN2FSuYihYqXZDrFmFTuds2EVUTiKIAgTUDREzMDBBHimDl2JWZUQBWZFyVAAARFahOT5N2uVxEEkCGh0/3qQI1VVWgMledWVWRVes9QgprCSMLuXrGXbQLdLrPMUWkUCFAoQTrXmJBIzMSGdFURERNfM6IkILHnHMi8/B8nFNgIppr7SNDIIGMhEKqIVInEJ4lEEkkuqAJMqVXzZkffPDxD37hq3/pAOCvfuGvfvbjd1WxVeGt53Yfj5/5LiebiYiIiOiHiwE0EREREX0ECvjDdz/77Tf3P/7cW4/XqJS3v/78H/zb3/vKe5//1tvvSPk2oiQt9quk5hSoR5WGVcmMBFRK1mRHrRnntYpcIlKSUgKt9U8lAoOJoQQKXbcLVZs1iEDU0ETFaw1pqApUUkXGuB7XI6usmbUWc0aVClai7eEoiEKbiqkAyCqRypKySkjK9DnmIaIlKMB6g9gMz6yI8BnIyLM13ZopKlUEJTj3MiLTRk6YwBOhjogqE4kqAFbm5U31MdQuc6D3q7Qa+STvvpVztwDm0Z+3F//9my//4IMP/uRPPtqnnYiIiIh+5jCAJiIiIqIfCwX87uff/tbbb/z+5z45e9cMC0lIFbISaxQZKZk94k0fH+BuWHatKYFYox5wgUAtI1pKWimqokQhqlIlkNJUIAVIUVWxFNWqFBFIAFUqkiKQTA8fx/V2vk8iEnlrGQNVmYi14CEC6CofA4D4KlHDI9JrXXCECLqaWmRUIlOg0IJa14BaWLZUdBUFEtf7F/rF3/rav/77n/1fn3wtK1HIrMxaOx8AUFIogUQBWq4CQAImaRGC6g/19P0//GieTiIiIiIiAAygiYiIiOgnzpff+/wj2hQZoqkJZKGkAJGVzMoaxDinN6rOw4a3/1bf34ledecCBJKCOt8MBFWZ4dPDM/J8y1VZCdT6q5BAldSZQQOAFIAECpWSWRmZWec7UxHT9aYyV19bVEShKqK3rWsViGTz/Ft//Ozt781f/tp3+SM7EREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREf04+D/5BQPQy/NfZwAAAABJRU5ErkJggg==" height="1080" preserveAspectRatio="xMidYMid meet"/></g></g></svg>
